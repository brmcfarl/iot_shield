//
// 
// PERMISSION IS HEREBY GRANTED, FREE OF CHARGE, TO ANY PERSON LEGALLY OBTAINING A COPY 
// OF THIS IP TO USE THE IP FOR THE PURPOSE OF THE DEVELOPMENT OF THE GALILEO CSI2 SHIELD,
// SUBJECT TO THE FOLLOWING CONDITIONS:
// 
// 1.	THE IP SHALL BE USED FOR THE PURPOSE STATED ABOVE, AND WILL NOT BE USED FOR ANY OTHER
// PURPOSE.
// 
// 2. THE USER WILL NOT REVERSE ENGINEER OR ATTEMPT TO REVERSE ENGINEER THE IP
// 
// 3. THE USER WILL NOT MODIFY OR OTHERWISE CREATE MODIFIED VERSIONS OF THE IP AND/OR OF
// PARTS THEREOF 
// 
// 4. THE FOLLOWING TEXT SHALL BE INCLUDED IN ALL COPIES OF THE IP:
// 
//                COPYRIGHT VLSI PLUS, LTD. 2014
// 
// 
// 5.	THE IP IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING 
// BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE 
// AND NONINFRINGEMENT. IN NO EVENT SHALL VLSI PLUS, LTD. BE LIABLE FOR ANY CLAIM, DAMAGES 
// OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, 
// OUT OF OR IN CONNECTION WITH THE IP OR THE USE OR OTHER DEALINGS IN THE IP.
//
//
////////////////////////////////////////////////////////////////////////////////////////////////////
//                              COPYRIGHT VLSI PLUS, LTD. 2014                                    //
////////////////////////////////////////////////////////////////////////////////////////////////////
// 9-April-2015 - two manual changes, plus version step-up (search for 9-April-2015)
module svr_lt2
(
svr_pixel,
svr_pixel_valid,
svr_channel_id,
svr_fs,
svr_fe,
svr_ls,
svr_le,
svr_data_type,
svr_cpu_int,
readdata,
fclk,
pclk,
reset_n,
address,
writedata,
write,
read,
lpck_p,
lpck_n,
lpd1_p,
lpd1_n,
hs_clk,
hs_d1,
hs_d2,
lpd2_p,
lpd2_n
);
output [9:0] svr_pixel;
output svr_pixel_valid;
output [1:0] svr_channel_id;
output svr_fs;
output svr_fe;
output svr_ls;
output svr_le;
output [5:0] svr_data_type;
output svr_cpu_int;
output [31:0] readdata;
input fclk;
input pclk;
input reset_n;
input [5:0] address;
input [31:0] writedata;
input write;
input read;
input lpck_p;
input lpck_n;
input lpd1_p;
input lpd1_n;
input hs_clk;
input hs_d1;
input hs_d2;
input lpd2_p;
input lpd2_n;

`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
// changed the version below (was 32'h01146101)
`define SVRJNvGI 			   32'h01154091
`define SVRHElWy 
`timescale 1ns/1ps

wire
[
7
:
0
]
SVRrpMRA
;
wire
[
7
:
0
]
SVRIhTvN
;
wire
SVRdxsDk
;
wire
SVRBlJoF
;
wire
SVRZyNzG
;
wire
SVRLFpfH
;
SVReJdvh
SVRCRBKD
(
.SVRaPJKf
(
pclk
)
,
.reset_n
(
reset_n
)
,
.SVRnXiwb
(
SVRZyNzG
)
,
.SVRSrADr
(
SVRLFpfH
)
)
;
wire
SVRWiNOI
,
SVRyEtuR
;
SVReJdvh
SVRmPjKv
(
.SVRaPJKf
(
pclk
)
,
.reset_n
(
reset_n
)
,
.SVRnXiwb
(
reset_n
)
,
.SVRSrADr
(
SVRWiNOI
)
)
;
SVReJdvh
SVRGUeSk
(
.SVRaPJKf
(
fclk
)
,
.reset_n
(
reset_n
)
,
.SVRnXiwb
(
reset_n
)
,
.SVRSrADr
(
SVRyEtuR
)
)
;
wire
SVRCqyoW
;
SVRAbIZo
SVRZTmsY
(
.SVRlqCbq
(
hs_clk
)
,
.SVRfiOaI
(
SVRZyNzG
)
,
.SVRoXPSh
(
hs_d1
)
,
.SVRHYuWd
(
SVRrpMRA
)
,
.SVRqzkYb
(
SVRdxsDk
)
)
;
SVRAbIZo
SVRImfZA
(
.SVRlqCbq
(
hs_clk
)
,
.SVRfiOaI
(
SVRCqyoW
)
,
.SVRoXPSh
(
hs_d2
)
,
.SVRHYuWd
(
SVRIhTvN
)
,
.SVRqzkYb
(
SVRBlJoF
)
)
;
wire
SVRrGCzn
=
(
write
|
read
)
;
wire
[
23
:
0
]
SVRujkFX
;
assign
svr_pixel
=
SVRujkFX
[
9
:
0
]
;
SVRWXaIp
SVRYyaRh
(
.svr_pixel
(
SVRujkFX
)
,
.svr_pixel_valid
(
svr_pixel_valid
)
,
.SVRgDTYn
(
svr_channel_id
)
,
.svr_fs
(
svr_fs
)
,
.svr_fe
(
svr_fe
)
,
.svr_ls
(
svr_ls
)
,
.svr_le
(
svr_le
)
,
.svr_data_type
(
svr_data_type
)
,
.svr_cpu_int
(
svr_cpu_int
)
,
.SVRTVbtZ
(
readdata
)
,
.SVRCqyoW
(
SVRCqyoW
)
,
.fclk
(
fclk
)
,
.pclk
(
pclk
)
,
.SVRrGCzn
(
SVRrGCzn
)
,
.SVRzMTVm
(
1'b1
)
,
.SVRWiNOI
(
SVRWiNOI
)
,
.SVRyEtuR
(
SVRyEtuR
)
,
.SVRyMsqX
(
address
)
,
.SVRmtjIy
(
writedata
)
,
.SVRSCAjD
(
write
)
,
.SVRIhjxF
(
lpck_p
)
,
.SVRdxaEg
(
lpck_n
)
,
.SVRBlapD
(
lpd1_p
)
,
.SVRZYVzf
(
lpd1_n
)
,
.SVRdxsDk
(
SVRdxsDk
)
,
.SVRrpMRA
(
SVRrpMRA
)
,
`ifdef SVRCadQw 
.SVRzZXMc
(
lpd2_p
)
,
.SVRYSUlS
(
lpd2_n
)
,
.SVRBlJoF
(
SVRBlJoF
)
,
.SVRIhTvN
(
SVRIhTvN
)
,
`endif
.SVRZyNzG
(
SVRZyNzG
)
)
;
endmodule
module SVRAbIZo
(
SVRlqCbq
,
SVRfiOaI
,
SVRoXPSh
,
SVRHYuWd
,
SVRqzkYb
)
;
input
SVRlqCbq
;
input
SVRfiOaI
;
input
SVRoXPSh
;
output
[
7
:
0
]
SVRHYuWd
;
output
SVRqzkYb
;
reg
[
3
:
0
]
SVRzwXfW
;
reg
[
3
:
0
]
SVRyEuVO
;
reg
[
7
:
0
]
SVRmpKxU
;
reg
[
1
:
0
]
SVRSaoeO
;
reg
SVRITCUK
,
SVRRwoxs
;
always
@
(
posedge
SVRlqCbq
)
SVRITCUK
<=
SVRoXPSh
;
always
@
(
negedge
SVRlqCbq
)
SVRRwoxs
<=
SVRoXPSh
;
wire
[
7
:
0
]
SVRHedea
=
SVRmpKxU
;
always
@
(
posedge
SVRlqCbq
or
negedge
SVRfiOaI
)
if
(
~SVRfiOaI
)
SVRSaoeO
[
1
:
0
]
<=
2'b00
;
else
SVRSaoeO
[
1
:
0
]
<=
SVRSaoeO
[
1
:
0
]
+
2'b01
;
always
@
(
posedge
SVRlqCbq
)
SVRyEuVO
[
3
:
0
]
<=
{
SVRITCUK
,
SVRyEuVO
[
3
:
1
]
}
;
always
@
(
negedge
SVRlqCbq
)
SVRzwXfW
[
3
:
0
]
<=
{
SVRRwoxs
,
SVRzwXfW
[
3
:
1
]
}
;
always
@
(
posedge
SVRlqCbq
)
begin
if
(
SVRSaoeO
[
1
:
0
]
==
2'b00
)
SVRmpKxU
[
7
:
0
]
<=
{
SVRzwXfW
[
3
]
,
SVRyEuVO
[
3
]
,
SVRzwXfW
[
2
]
,
SVRyEuVO
[
2
]
,
SVRzwXfW
[
1
]
,
SVRyEuVO
[
1
]
,
SVRzwXfW
[
0
]
,
SVRyEuVO
[
0
]
}
;
else
SVRmpKxU
[
7
:
0
]
<=
SVRHedea
[
7
:
0
]
;
end
assign
SVRqzkYb
=
SVRSaoeO
[
1
]
;
reg
[
7
:
0
]
SVRHYuWd
;
initial
#
0
SVRHYuWd
=
8'd0
;
always
@
(
posedge
SVRlqCbq
)
SVRHYuWd
<=
SVRHedea
;
endmodule
module SVReJdvh
(
SVRaPJKf
,
reset_n
,
SVRnXiwb
,
SVRSrADr
)
;
input
SVRaPJKf
,
reset_n
,
SVRnXiwb
;
output
SVRSrADr
;
reg
[
1
:
0
]
SVRCvxUQ
;
always
@
(
posedge
SVRaPJKf
or
negedge
reset_n
)
if
(
~reset_n
)
SVRCvxUQ
<=
2'b00
;
else
SVRCvxUQ
<=
{
SVRCvxUQ
[
0
]
,
SVRnXiwb
}
;
assign
SVRSrADr
=
SVRCvxUQ
[
1
]
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRWXaIp
(
svr_pixel
,
svr_pixel_valid
,
SVRgDTYn
,
svr_fs
,
svr_fe
,
svr_ls
,
svr_le
,
svr_data_type
,
svr_cpu_int
,
SVRTVbtZ
,
SVRCqyoW
,
fclk
,
pclk
,
SVRrGCzn
,
SVRzMTVm
,
SVRWiNOI
,
SVRyEtuR
,
SVRyMsqX
,
SVRmtjIy
,
SVRSCAjD
,
SVRIhjxF
,
SVRdxaEg
,
SVRBlapD
,
SVRZYVzf
,
SVRdxsDk
,
SVRrpMRA
,
SVRzZXMc
,
SVRYSUlS
,
SVRBlJoF
,
SVRIhTvN
,
SVRZyNzG
)
;
output
[
23
:
0
]
svr_pixel
;
output
svr_pixel_valid
;
output
[
1
:
0
]
SVRgDTYn
;
output
svr_fs
;
output
svr_fe
;
output
svr_ls
;
output
svr_le
;
output
[
5
:
0
]
svr_data_type
;
output
svr_cpu_int
;
output
[
31
:
0
]
SVRTVbtZ
;
output
SVRCqyoW
;
input
fclk
;
input
pclk
;
input
SVRrGCzn
;
input
SVRzMTVm
;
input
SVRWiNOI
;
input
SVRyEtuR
;
input
[
5
:
0
]
SVRyMsqX
;
input
[
31
:
0
]
SVRmtjIy
;
input
SVRSCAjD
;
input
SVRIhjxF
;
input
SVRdxaEg
;
input
SVRBlapD
;
input
SVRZYVzf
;
input
SVRdxsDk
;
input
[
7
:
0
]
SVRrpMRA
;
input
SVRzZXMc
;
input
SVRYSUlS
;
input
SVRBlJoF
;
input
[
7
:
0
]
SVRIhTvN
;
output
SVRZyNzG
;
wire
[
7
:
0
]
SVRfxZHB
;
wire
SVROEvJE
;
wire
SVRuPKrP
;
wire
SVRWnoBL
;
wire
SVRYgHNS
;
wire
SVRLwmmN
;
wire
SVRslgGT
;
wire
SVRVYyIN
;
wire
SVRJsIJK
;
wire
[
7
:
0
]
SVRrjRrs
;
wire
SVRUxrba
;
wire
SVRjFeTQ
;
wire
SVRQiYom
;
wire
[
27
:
0
]
SVRHXUZw
;
wire
SVRcstsC
;
wire
SVRnCFbF
;
wire
SVRgOPAP
;
wire
SVRdUuNu
;
wire
SVRbxKtK
;
wire
SVRAlSjs
;
wire
SVRNfWej
;
wire
SVRTcyCe
;
SVRIUHgT
SVRDQMvn
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRIhjxF
)
,
.SVRnHHOy
(
SVRgOPAP
)
)
;
SVRIUHgT
SVRSJMmd
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRdxaEg
)
,
.SVRnHHOy
(
SVRdUuNu
)
)
;
SVRIUHgT
SVRilPyS
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRBlapD
)
,
.SVRnHHOy
(
SVRbxKtK
)
)
;
SVRIUHgT
SVREFumw
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRZYVzf
)
,
.SVRnHHOy
(
SVRAlSjs
)
)
;
SVRIUHgT
SVRbjGYb
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRzZXMc
)
,
.SVRnHHOy
(
SVRNfWej
)
)
;
SVRIUHgT
SVRMXLRR
(
.SVRaPJKf
(
fclk
)
,
.SVRAopDX
(
SVRYSUlS
)
,
.SVRnHHOy
(
SVRTcyCe
)
)
;
wire
SVRfSoOm
;
wire
SVRopDmx
;
wire
SVRTAKyC
;
wire
SVRIgOeF
;
SVRDWPuG
SVRoYukQ
(
.SVRcstsC
(
SVRcstsC
)
,
.SVRZyNzG
(
SVRZyNzG
)
,
.SVRfSoOm
(
SVRfSoOm
)
,
.fclk
(
fclk
)
,
.pclk
(
pclk
)
,
.SVRrGCzn
(
SVRrGCzn
)
,
.SVRzMTVm
(
SVRzMTVm
)
,
.SVRWiNOI
(
SVRWiNOI
)
,
.SVRyEtuR
(
SVRyEtuR
)
,
.SVRyMsqX
(
SVRyMsqX
)
,
.SVRmtjIy
(
SVRmtjIy
[
31
:
0
]
)
,
.SVRSCAjD
(
SVRSCAjD
)
,
.SVRhzkfv
(
SVRfxZHB
[
7
:
0
]
)
,
.SVRuPKrP
(
SVRuPKrP
)
,
.SVRYgHNS
(
SVRYgHNS
)
,
.SVRWnoBL
(
SVRWnoBL
)
,
.SVRLwmmN
(
SVRLwmmN
)
,
.SVRVYyIN
(
SVRVYyIN
)
,
.SVRJsIJK
(
SVRJsIJK
)
,
.SVRopDmx
(
SVRopDmx
)
,
.SVROEvJE
(
SVROEvJE
)
,
.SVRnCFbF
(
SVRnCFbF
)
,
.svr_pixel
(
svr_pixel
[
23
:
0
]
)
,
.svr_pixel_valid
(
svr_pixel_valid
)
,
.SVRgDTYn
(
SVRgDTYn
)
,
.svr_fs
(
svr_fs
)
,
.svr_fe
(
svr_fe
)
,
.svr_ls
(
svr_ls
)
,
.svr_le
(
svr_le
)
,
.svr_data_type
(
svr_data_type
[
5
:
0
]
)
,
.svr_cpu_int
(
svr_cpu_int
)
,
.SVRTVbtZ
(
SVRTVbtZ
[
31
:
0
]
)
,
.SVRHXUZw
(
SVRHXUZw
[
27
:
0
]
)
,
.SVRCqyoW
(
SVRCqyoW
)
,
.SVRDmFCK
(
SVRrjRrs
[
7
:
0
]
)
,
.SVRjFeTQ
(
SVRjFeTQ
)
,
.SVRIgOeF
(
SVRIgOeF
)
,
.SVRQiYom
(
SVRQiYom
)
,
.SVRTAKyC
(
SVRTAKyC
)
,
.SVRUxrba
(
SVRUxrba
)
)
;
assign
SVRcstsC
=
~SVRZyNzG
;
SVRoGpos
SVRtJDZZ
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRZyNzG
(
SVRZyNzG
)
,
.SVRCqyoW
(
SVRCqyoW
)
,
.SVRfSoOm
(
SVRfSoOm
)
,
.SVRIhjxF
(
SVRgOPAP
)
,
.SVRdxaEg
(
SVRdUuNu
)
,
.SVRBlapD
(
SVRbxKtK
)
,
.SVRZYVzf
(
SVRAlSjs
)
,
.SVRdxsDk
(
SVRdxsDk
)
,
.SVRrpMRA
(
SVRrpMRA
[
7
:
0
]
)
,
.SVRHXUZw
(
SVRHXUZw
)
,
.SVRfxZHB
(
SVRfxZHB
[
7
:
0
]
)
,
.SVRRvUZM
(
SVRuPKrP
)
,
.SVRYgHNS
(
SVRYgHNS
)
,
.SVRWnoBL
(
SVRWnoBL
)
,
.SVRVYyIN
(
SVRVYyIN
)
,
.SVRJsIJK
(
SVRJsIJK
)
,
.SVRopDmx
(
SVRopDmx
)
,
.SVROEvJE
(
SVROEvJE
)
,
.SVRnCFbF
(
SVRnCFbF
)
,
.SVRLwmmN
(
SVRLwmmN
)
,
.SVRzZXMc
(
SVRNfWej
)
,
.SVRYSUlS
(
SVRTcyCe
)
,
.SVRBlJoF
(
SVRBlJoF
)
,
.SVRIhTvN
(
SVRIhTvN
[
7
:
0
]
)
,
.SVRrjRrs
(
SVRrjRrs
[
7
:
0
]
)
,
.SVRVkXzt
(
SVRjFeTQ
)
,
.SVRIgOeF
(
SVRIgOeF
)
,
.SVRQiYom
(
SVRQiYom
)
,
.SVRTAKyC
(
SVRTAKyC
)
,
.SVRUxrba
(
SVRUxrba
)
,
.SVRslgGT
(
SVRslgGT
)
)
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRIUHgT
(
SVRaPJKf
,
SVRAopDX
,
SVRnHHOy
)
;
input
SVRaPJKf
;
input
SVRAopDX
;
output
SVRnHHOy
;
reg
SVRVoBcb
;
wire
SVRJAJtr
,
SVRrNRJI
,
SVRITVrr
;
SVRRWXII
SVRvYyrr
(
.SVRSrADr
(
SVRJAJtr
)
,
.SVRnXiwb
(
SVRAopDX
)
,
.SVRlqCbq
(
SVRaPJKf
)
)
;
SVRRWXII
SVRkzMIi
(
.SVRSrADr
(
SVRrNRJI
)
,
.SVRnXiwb
(
SVRJAJtr
)
,
.SVRlqCbq
(
SVRaPJKf
)
)
;
SVRRWXII
SVRRfPjV
(
.SVRSrADr
(
SVRITVrr
)
,
.SVRnXiwb
(
SVRrNRJI
)
,
.SVRlqCbq
(
SVRaPJKf
)
)
;
wire
[
2
:
0
]
SVRVCUEx
=
{
SVRITVrr
,
SVRrNRJI
,
SVRJAJtr
}
;
initial
#
0
SVRVoBcb
=
1'b0
;
always
@
(
posedge
SVRaPJKf
)
`ifdef SVRxoxPL 
if
(
(
SVRVCUEx
==
3'b111
)
===
1'bx
)
SVRVoBcb
<=
1'bx
;
else
`endif
if
(
SVRVCUEx
==
3'b111
)
SVRVoBcb
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
SVRVCUEx
==
3'b000
)
===
1'bx
)
SVRVoBcb
<=
1'bx
;
`endif
else
if
(
SVRVCUEx
==
3'b000
)
SVRVoBcb
<=
1'b0
;
assign
SVRnHHOy
=
SVRVoBcb
;
endmodule
module SVRRWXII
(
SVRSrADr
,
SVRnXiwb
,
SVRlqCbq
)
;
output
reg
SVRSrADr
;
input
SVRnXiwb
,
SVRlqCbq
;
initial
SVRSrADr
=
1'b0
;
always
@
(
posedge
SVRlqCbq
)
SVRSrADr
<=
SVRnXiwb
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRoGpos
(
fclk
,
SVRJROZz
,
SVRZyNzG
,
SVRCqyoW
,
SVRfSoOm
,
SVRIhjxF
,
SVRdxaEg
,
SVRBlapD
,
SVRZYVzf
,
SVRdxsDk
,
SVRrpMRA
,
SVRHXUZw
,
SVRfxZHB
,
SVRRvUZM
,
SVRYgHNS
,
SVRWnoBL
,
SVRVYyIN
,
SVRJsIJK
,
SVRopDmx
,
SVROEvJE
,
SVRnCFbF
,
SVRLwmmN
,
SVRzZXMc
,
SVRYSUlS
,
SVRBlJoF
,
SVRIhTvN
,
SVRrjRrs
,
SVRVkXzt
,
SVRIgOeF
,
SVRQiYom
,
SVRTAKyC
,
SVRUxrba
,
SVRslgGT
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRZyNzG
;
input
SVRCqyoW
;
input
SVRfSoOm
;
input
SVRIhjxF
;
input
SVRdxaEg
;
input
SVRBlapD
;
input
SVRZYVzf
;
input
SVRdxsDk
;
input
[
7
:
0
]
SVRrpMRA
;
input
[
27
:
0
]
SVRHXUZw
;
output
[
7
:
0
]
SVRfxZHB
;
output
SVRRvUZM
;
output
SVRYgHNS
;
output
SVRWnoBL
;
output
SVRVYyIN
;
output
SVRJsIJK
;
output
SVRopDmx
;
output
SVROEvJE
;
output
SVRnCFbF
;
output
SVRLwmmN
;
input
SVRzZXMc
;
input
SVRYSUlS
;
input
SVRBlJoF
;
input
[
7
:
0
]
SVRIhTvN
;
output
[
7
:
0
]
SVRrjRrs
;
output
SVRVkXzt
;
output
SVRIgOeF
;
output
SVRQiYom
;
output
SVRTAKyC
;
output
SVRUxrba
;
output
SVRslgGT
;
wire
SVRLljSa
=
SVRZyNzG
;
wire
SVRezAor
=
SVRZyNzG
;
reg
[
2
:
0
]
SVROfJzz
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVROfJzz
<=
3'b000
;
else
if
(
SVRZyNzG
==
1'b0
)
SVROfJzz
<=
3'b000
;
else
if
(
SVRezAor
==
1'b0
)
SVROfJzz
<=
3'b000
;
else
SVROfJzz
<=
{
SVROfJzz
[
1
:
0
]
,
1'b1
}
;
wire
SVRgwnFd
=
SVROfJzz
[
2
]
;
wire
[
5
:
0
]
SVRpEcIs
;
wire
SVRtixjA
=
SVRIhjxF
;
wire
SVRvxhXD
=
SVRdxaEg
;
wire
SVRcstsC
=
~SVRZyNzG
;
SVRWEZQF
SVRKIVNG
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRcstsC
(
SVRcstsC
)
,
.SVRfiOaI
(
SVRLljSa
)
,
.SVREKtmH
(
SVRBlapD
)
,
.SVRBLFyH
(
SVRZYVzf
)
,
.SVRNSpMQ
(
SVRdxsDk
)
,
.SVRFPDlm
(
SVRrpMRA
)
,
.SVRHXUZw
(
SVRHXUZw
)
,
.SVRpEcIs
(
SVRpEcIs
)
,
.SVRbOkYW
(
SVRfxZHB
)
,
.SVRmnBrp
(
SVRRvUZM
)
,
.SVRGGNIH
(
SVRYgHNS
)
,
.SVRqQtRq
(
SVRJsIJK
)
,
.SVRuOfoz
(
SVRopDmx
)
,
.SVRkUcHM
(
SVROEvJE
)
,
.SVRfxBqT
(
SVRLwmmN
)
)
;
SVRWEZQF
SVROEJAn
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRcstsC
(
SVRcstsC
)
,
.SVRfiOaI
(
SVRCqyoW
)
,
.SVREKtmH
(
SVRzZXMc
)
,
.SVRBLFyH
(
SVRYSUlS
)
,
.SVRNSpMQ
(
SVRBlJoF
)
,
.SVRFPDlm
(
SVRIhTvN
)
,
.SVRHXUZw
(
SVRHXUZw
)
,
.SVRpEcIs
(
SVRpEcIs
)
,
.SVRbOkYW
(
SVRrjRrs
)
,
.SVRmnBrp
(
SVRVkXzt
)
,
.SVRGGNIH
(
SVRIgOeF
)
,
.SVRqQtRq
(
SVRQiYom
)
,
.SVRuOfoz
(
SVRTAKyC
)
,
.SVRkUcHM
(
SVRUxrba
)
,
.SVRfxBqT
(
SVRslgGT
)
)
;
SVRuPrNG
SVRuPrNG
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRcstsC
(
SVRcstsC
)
,
.SVRfiOaI
(
SVRgwnFd
)
,
.SVRWNemH
(
SVRtixjA
)
,
.SVRknyyH
(
SVRvxhXD
)
,
.SVRRZHEh
(
SVRHXUZw
[
23
:
16
]
)
,
.SVRGGNIH
(
SVRWnoBL
)
,
.SVRhTMHu
(
SVRVYyIN
)
)
;
wire
SVRDwTqK
;
SVRAESaj
SVRnpwAe
(
.SVRnXiwb
(
SVRdxsDk
)
,
.SVRlqCbq
(
fclk
)
,
.SVRGhlnc
(
SVRDwTqK
)
)
;
reg
[
5
:
0
]
SVRcxbZr
,
SVRNEWRz
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRcxbZr
<=
6'b000000
;
else
if
(
SVRcstsC
==
1'b1
)
SVRcxbZr
<=
6'b000000
;
else
if
(
SVRRvUZM
)
SVRcxbZr
<=
6'b000000
;
else
SVRcxbZr
<=
SVRcxbZr
+
6'b000001
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRNEWRz
<=
6'b000000
;
else
if
(
SVRcstsC
==
1'b1
)
SVRNEWRz
<=
6'b000000
;
else
if
(
SVRRvUZM
)
SVRNEWRz
<=
SVRcxbZr
;
assign
SVRpEcIs
=
SVRNEWRz
;
wire
SVRtpYVm
;
SVRAESaj
SVRJhZxg
(
.SVRnXiwb
(
~SVRdxsDk
)
,
.SVRlqCbq
(
fclk
)
,
.SVRGhlnc
(
SVRtpYVm
)
)
;
wire
SVRRDZlD
=
SVRDwTqK
|
SVRtpYVm
;
wire
SVRnCFbF
;
reg
[
4
:
0
]
SVRVOZFo
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRVOZFo
<=
5'b00000
;
else
if
(
SVRcstsC
==
1'b1
)
SVRVOZFo
<=
5'b00000
;
else
if
(
(
SVRfSoOm
==
1'b1
)
&&
(
SVRYgHNS
==
1'b0
)
)
SVRVOZFo
<=
5'b00000
;
else
if
(
SVRgwnFd
)
begin
if
(
SVRRDZlD
)
SVRVOZFo
<=
5'b00000
;
else
SVRVOZFo
<=
SVRVOZFo
+
5'b00001
;
end
else
SVRVOZFo
<=
5'b00000
;
assign
SVRnCFbF
=
SVRgwnFd
&
(
SVRVOZFo
==
{
SVRHXUZw
[
27
:
24
]
,
1'b0
}
)
;
endmodule
module SVRAESaj
(
SVRnXiwb
,
SVRlqCbq
,
SVRGhlnc
)
;
input
SVRnXiwb
;
input
SVRlqCbq
;
output
SVRGhlnc
;
reg
SVRxUZph
;
wire
SVRlXZHd
;
reg
SVRFYZQb
;
initial
#
0
SVRxUZph
=
1'b0
;
always
@
(
posedge
SVRnXiwb
)
SVRxUZph
<=
~SVRxUZph
;
SVRBSVNR
SVRnWXTv
(
.SVRgYYWK
(
SVRxUZph
)
,
.SVRpsVqj
(
SVRlqCbq
)
,
.SVRtCTAv
(
SVRlXZHd
)
)
;
initial
#
0
SVRFYZQb
=
1'b0
;
always
@
(
posedge
SVRlqCbq
)
SVRFYZQb
<=
SVRlXZHd
;
assign
SVRGhlnc
=
SVRlXZHd
^
SVRFYZQb
;
endmodule
module SVRvHSFb
(
SVRKqWPA
,
SVRgYYWK
,
SVRtCTAv
,
SVRpsVqj
)
;
input
SVRKqWPA
;
input
SVRgYYWK
;
input
SVRpsVqj
;
output
SVRtCTAv
;
reg
SVRsiYun
;
reg
SVRtCTAv
;
always
@
(
posedge
SVRpsVqj
or
posedge
SVRKqWPA
)
if
(
SVRKqWPA
)
begin
SVRsiYun
<=
1'b0
;
SVRtCTAv
<=
1'b0
;
end
else
begin
SVRsiYun
<=
SVRgYYWK
;
SVRtCTAv
<=
SVRsiYun
;
end
endmodule
module SVRWEZQF
(
fclk
,
SVRJROZz
,
SVRcstsC
,
SVRfiOaI
,
SVREKtmH
,
SVRBLFyH
,
SVRNSpMQ
,
SVRFPDlm
,
SVRHXUZw
,
SVRpEcIs
,
SVRbOkYW
,
SVRmnBrp
,
SVRGGNIH
,
SVRqQtRq
,
SVRuOfoz
,
SVRkUcHM
,
SVRfxBqT
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRcstsC
;
input
SVRfiOaI
;
input
SVREKtmH
;
input
SVRBLFyH
;
input
SVRNSpMQ
;
input
[
7
:
0
]
SVRFPDlm
;
input
[
27
:
0
]
SVRHXUZw
;
input
[
5
:
0
]
SVRpEcIs
;
output
[
7
:
0
]
SVRbOkYW
;
output
SVRmnBrp
;
output
SVRGGNIH
;
output
SVRqQtRq
;
output
SVRuOfoz
;
output
SVRkUcHM
;
output
SVRfxBqT
;
reg
[
2
:
0
]
SVRjezKG
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRjezKG
<=
3'b000
;
else
if
(
SVRcstsC
==
1'b1
)
SVRjezKG
<=
3'b000
;
else
if
(
SVRfiOaI
==
1'b0
)
SVRjezKG
<=
3'b000
;
else
SVRjezKG
<=
{
SVRjezKG
[
1
:
0
]
,
1'b1
}
;
wire
SVReCmsq
=
SVRjezKG
[
2
]
;
wire
SVRuOfoz
;
wire
SVRcogji
;
wire
SVRWNemH
=
SVREKtmH
;
wire
SVRknyyH
=
SVRBLFyH
;
wire
SVRnaZWU
;
wire
SVRgAzyx
;
wire
[
7
:
0
]
SVRpGIEC
;
wire
SVRhqrpO
;
SVRpBeaL
SVRpBeaL
(
.SVRJROZz
(
SVRJROZz
)
,
.SVRHncAS
(
SVRNSpMQ
)
,
.SVRcaxfN
(
SVRFPDlm
)
,
.write
(
SVRfiOaI
)
,
.SVRaNsOW
(
fclk
)
,
.SVRMmFmp
(
SVRpGIEC
)
,
.SVRhqrpO
(
SVRhqrpO
)
)
;
wire
SVRtGpGH
,
SVRvJDIH
,
SVRWKKJH
,
SVRysSRq
,
SVRmjWvi
,
SVRGeYkE
,
SVRqczfp
,
SVRuuivY
;
wire
SVRkkEkz
,
SVRffpFM
,
SVRCCHpt
,
SVRAHmAa
,
SVRZjCfr
,
SVRlYjvZ
,
SVRrSaDq
,
SVRupWgz
;
reg
[
6
:
0
]
SVRKhyDM
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
~SVRJROZz
)
SVRKhyDM
<=
7'd0
;
else
if
(
SVRhqrpO
)
SVRKhyDM
<=
SVRpGIEC
[
7
:
1
]
;
wire
[
14
:
0
]
SVRSdMot
=
{
SVRpGIEC
,
SVRKhyDM
}
;
SVRiVOzA
SVRExUmN
(
.SVRbfTyK
(
SVRSdMot
[
14
:
7
]
)
,
.SVRMvSeJ
(
SVRtGpGH
)
,
.SVRfeSui
(
SVRkkEkz
)
)
;
SVRiVOzA
SVRoVRcv
(
.SVRbfTyK
(
SVRSdMot
[
13
:
6
]
)
,
.SVRMvSeJ
(
SVRvJDIH
)
,
.SVRfeSui
(
SVRffpFM
)
)
;
SVRiVOzA
SVRTQRtB
(
.SVRbfTyK
(
SVRSdMot
[
12
:
5
]
)
,
.SVRMvSeJ
(
SVRWKKJH
)
,
.SVRfeSui
(
SVRCCHpt
)
)
;
SVRiVOzA
SVRIOrCE
(
.SVRbfTyK
(
SVRSdMot
[
11
:
4
]
)
,
.SVRMvSeJ
(
SVRysSRq
)
,
.SVRfeSui
(
SVRAHmAa
)
)
;
SVRiVOzA
SVRrUioP
(
.SVRbfTyK
(
SVRSdMot
[
10
:
3
]
)
,
.SVRMvSeJ
(
SVRmjWvi
)
,
.SVRfeSui
(
SVRZjCfr
)
)
;
SVRiVOzA
SVRixeHu
(
.SVRbfTyK
(
SVRSdMot
[
9
:
2
]
)
,
.SVRMvSeJ
(
SVRGeYkE
)
,
.SVRfeSui
(
SVRlYjvZ
)
)
;
SVRiVOzA
SVRElCqK
(
.SVRbfTyK
(
SVRSdMot
[
8
:
1
]
)
,
.SVRMvSeJ
(
SVRqczfp
)
,
.SVRfeSui
(
SVRrSaDq
)
)
;
SVRiVOzA
SVRbZJaj
(
.SVRbfTyK
(
SVRSdMot
[
7
:
0
]
)
,
.SVRMvSeJ
(
SVRuuivY
)
,
.SVRfeSui
(
SVRupWgz
)
)
;
wire
[
7
:
0
]
SVRAZrAE
=
{
SVRuuivY
,
SVRqczfp
,
SVRGeYkE
,
SVRmjWvi
,
SVRysSRq
,
SVRWKKJH
,
SVRvJDIH
,
SVRtGpGH
}
;
wire
[
7
:
0
]
SVRNZinP
=
{
SVRupWgz
,
SVRrSaDq
,
SVRlYjvZ
,
SVRZjCfr
,
SVRAHmAa
,
SVRCCHpt
,
SVRffpFM
,
SVRkkEkz
}
;
wire
[
2
:
0
]
SVRftazl
;
assign
SVRftazl
=
(
SVRAZrAE
[
7
]
)
?
3'd7
:
(
SVRAZrAE
[
6
]
)
?
3'd6
:
(
SVRAZrAE
[
5
]
)
?
3'd5
:
(
SVRAZrAE
[
4
]
)
?
3'd4
:
(
SVRAZrAE
[
3
]
)
?
3'd3
:
(
SVRAZrAE
[
2
]
)
?
3'd2
:
(
SVRAZrAE
[
1
]
)
?
3'd1
:
(
SVRAZrAE
[
0
]
)
?
3'd0
:
3'd0
;
reg
[
2
:
0
]
SVROcWEw
;
reg
[
2
:
0
]
SVRubypl
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRubypl
<=
3'b000
;
else
if
(
SVRcstsC
)
SVRubypl
<=
3'b000
;
else
if
(
(
(
|
SVRAZrAE
)
&&
SVRcogji
&&
(
SVROcWEw
==
3'b000
)
)
)
SVRubypl
<=
SVRftazl
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVROcWEw
<=
3'b000
;
else
if
(
SVRcstsC
==
1'b1
)
SVROcWEw
<=
3'b000
;
else
if
(
SVRqQtRq
)
SVROcWEw
<=
3'b000
;
else
if
(
(
~
(
|
SVRAZrAE
)
|
~SVRcogji
)
&&
(
SVROcWEw
==
3'b000
)
)
SVROcWEw
<=
3'b000
;
else
if
(
(
|
(
SVRAZrAE
&
(
~SVRNZinP
)
)
)
&&
SVRcogji
&&
(
SVROcWEw
==
3'b000
)
&&
SVRhqrpO
)
SVROcWEw
<=
3'b011
;
else
if
(
(
|
(
SVRNZinP
&
SVRAZrAE
)
)
&&
SVRcogji
&&
(
SVROcWEw
==
3'b000
)
&&
SVRhqrpO
)
SVROcWEw
<=
3'b111
;
else
if
(
(
SVROcWEw
[
1
:
0
]
==
2'b11
)
)
SVROcWEw
<=
3'b001
;
assign
SVRfxBqT
=
(
SVROcWEw
[
1
:
0
]
==
2'b11
)
?
1'b1
:
1'b0
;
assign
SVRuOfoz
=
(
SVROcWEw
==
3'b111
)
?
1'b1
:
1'b0
;
wire
[
7
:
0
]
SVRWThAW
;
assign
SVRWThAW
=
(
SVRnaZWU
==
1'b0
)
?
8'h00
:
(
SVRubypl
[
2
:
0
]
==
3'b000
)
?
SVRSdMot
[
14
:
7
]
:
(
SVRubypl
[
2
:
0
]
==
3'b001
)
?
SVRSdMot
[
13
:
6
]
:
(
SVRubypl
[
2
:
0
]
==
3'b010
)
?
SVRSdMot
[
12
:
5
]
:
(
SVRubypl
[
2
:
0
]
==
3'b011
)
?
SVRSdMot
[
11
:
4
]
:
(
SVRubypl
[
2
:
0
]
==
3'b100
)
?
SVRSdMot
[
10
:
3
]
:
(
SVRubypl
[
2
:
0
]
==
3'b101
)
?
SVRSdMot
[
9
:
2
]
:
(
SVRubypl
[
2
:
0
]
==
3'b110
)
?
SVRSdMot
[
8
:
1
]
:
(
SVRubypl
[
2
:
0
]
==
3'b111
)
?
SVRSdMot
[
7
:
0
]
:
SVRSdMot
[
7
:
0
]
;
reg
[
7
:
0
]
SVRbOkYW
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
~SVRJROZz
)
SVRbOkYW
<=
8'd0
;
else
if
(
SVRhqrpO
)
SVRbOkYW
<=
SVRWThAW
;
reg
SVRYWdnY
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
~SVRJROZz
)
SVRYWdnY
<=
1'b0
;
else
SVRYWdnY
<=
SVRhqrpO
;
assign
SVRmnBrp
=
(
SVRfxBqT
)
?
1'b0
:
(
SVRgAzyx
==
1'b0
)
?
1'b0
:
SVRYWdnY
;
SVRzYBgZ
SVRzYBgZ
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRcstsC
(
SVRcstsC
)
,
.SVRfiOaI
(
SVReCmsq
)
,
.SVRWNemH
(
SVRWNemH
)
,
.SVRknyyH
(
SVRknyyH
)
,
.SVRRZHEh
(
SVRHXUZw
[
15
:
8
]
)
,
.SVRySJvq
(
SVRfxBqT
)
,
.SVRpEcIs
(
SVRpEcIs
[
5
:
0
]
)
,
.SVRgAzyx
(
SVRgAzyx
)
,
.SVRcogji
(
SVRcogji
)
,
.SVRGGNIH
(
SVRGGNIH
)
,
.SVRhTMHu
(
SVRqQtRq
)
,
.SVRnaZWU
(
SVRnaZWU
)
,
.SVRfeSui
(
SVRkUcHM
)
)
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRiVOzA
(
SVRbfTyK
,
SVRMvSeJ
,
SVRfeSui
`ifdef SVRsQYvh 
,
SVRvovDu
`endif
)
;
input
wire
[
7
:
0
]
SVRbfTyK
;
output
SVRMvSeJ
;
output
SVRfeSui
;
`ifdef SVRsQYvh 
input
wire
[
7
:
0
]
SVRvovDu
;
`endif
`ifdef SVRsQYvh 
wire
[
7
:
0
]
SVRkHKoK
=
SVRbfTyK
^
SVRvovDu
;
`else
wire
[
7
:
0
]
SVRkHKoK
=
{
~SVRbfTyK
[
7
]
,
SVRbfTyK
[
6
]
,
~SVRbfTyK
[
5
]
,
~SVRbfTyK
[
4
]
,
~SVRbfTyK
[
3
]
,
SVRbfTyK
[
2
]
,
SVRbfTyK
[
1
]
,
SVRbfTyK
[
0
]
}
;
`endif
wire
[
1
:
0
]
SVRRjOZI
=
{
1'b0
,
SVRkHKoK
[
0
]
}
+
{
1'b0
,
SVRkHKoK
[
1
]
}
;
wire
[
1
:
0
]
SVRVeUzR
=
{
1'b0
,
SVRkHKoK
[
2
]
}
+
{
1'b0
,
SVRkHKoK
[
3
]
}
+
{
1'b0
,
SVRkHKoK
[
4
]
}
;
wire
[
1
:
0
]
SVRxcXMV
=
{
1'b0
,
SVRkHKoK
[
5
]
}
+
{
1'b0
,
SVRkHKoK
[
6
]
}
+
{
1'b0
,
SVRkHKoK
[
7
]
}
;
wire
[
3
:
0
]
SVRlByTx
=
{
2'b00
,
SVRRjOZI
}
+
{
2'b00
,
SVRVeUzR
}
+
{
2'b00
,
SVRxcXMV
}
;
assign
SVRMvSeJ
=
(
SVRlByTx
[
3
:
1
]
==
3'd0
)
?
1'b1
:
1'b0
;
assign
SVRfeSui
=
(
SVRlByTx
!=
4'd0
)
?
1'b1
:
1'b0
;
endmodule
module SVRpBeaL
(
SVRJROZz
,
SVRHncAS
,
SVRcaxfN
,
write
,
SVRaNsOW
,
SVRMmFmp
,
SVRhqrpO
)
;
input
SVRJROZz
;
input
SVRHncAS
;
input
[
7
:
0
]
SVRcaxfN
;
input
write
;
input
SVRaNsOW
;
output
[
7
:
0
]
SVRMmFmp
;
output
SVRhqrpO
;
reg
[
7
:
0
]
SVRMmFmp
;
reg
SVRhqrpO
;
wire
SVRRgiPc
,
SVRHWZms
;
assign
SVRHWZms
=
~SVRRgiPc
;
wire
[
7
:
0
]
SVRpGIEC
;
SVRCRVYZ
#
8
SVRaPTRq
(
.reset_n
(
SVRJROZz
)
,
.SVRHncAS
(
SVRHncAS
)
,
.SVRAUWvI
(
SVRcaxfN
)
,
.SVRnxYkr
(
write
)
,
.SVRaNsOW
(
SVRaNsOW
)
,
.SVRGlzFI
(
SVRHWZms
)
,
.SVRcziii
(
SVRpGIEC
)
,
.SVRRgiPc
(
SVRRgiPc
)
)
;
always
@
(
posedge
SVRaNsOW
)
SVRMmFmp
<=
SVRpGIEC
;
always
@
(
posedge
SVRaNsOW
)
SVRhqrpO
<=
~SVRRgiPc
;
endmodule
module SVRCRVYZ
(
reset_n
,
SVRHncAS
,
SVRAUWvI
,
SVRnxYkr
,
SVRaNsOW
,
SVRGlzFI
,
SVRcziii
,
SVRRgiPc
)
;
parameter
SVRBmeeE
=
32
;
input
reset_n
;
input
SVRHncAS
;
input
[
SVRBmeeE
-
1
:
0
]
SVRAUWvI
;
input
SVRnxYkr
;
input
SVRaNsOW
;
input
SVRGlzFI
;
output
[
SVRBmeeE
-
1
:
0
]
SVRcziii
;
output
SVRRgiPc
;
reg
[
SVRBmeeE
-
1
:
0
]
SVRngccP
[
7
:
0
]
;
reg
[
3
:
0
]
SVRsWwtl
;
always
@
(
posedge
SVRHncAS
or
negedge
reset_n
)
if
(
~reset_n
)
SVRsWwtl
<=
4'd0
;
else
if
(
SVRnxYkr
)
SVRsWwtl
<=
SVRsWwtl
+
4'd1
;
reg
[
3
:
0
]
SVRjyLJF
;
always
@
(
posedge
SVRaNsOW
or
negedge
reset_n
)
if
(
~reset_n
)
SVRjyLJF
<=
4'd0
;
else
if
(
(
SVRGlzFI
)
&&
(
~SVRRgiPc
)
)
SVRjyLJF
<=
SVRjyLJF
+
4'd1
;
always
@
(
posedge
SVRHncAS
)
if
(
SVRnxYkr
)
SVRngccP
[
SVRsWwtl
[
2
:
0
]
]
<=
SVRAUWvI
;
assign
SVRcziii
=
SVRngccP
[
SVRjyLJF
[
2
:
0
]
]
;
wire
[
3
:
0
]
SVReMSRP
=
(
SVRsWwtl
==
4'b0000
)
?
4'b0000
:
(
SVRsWwtl
==
4'b0001
)
?
4'b0001
:
(
SVRsWwtl
==
4'b0010
)
?
4'b0011
:
(
SVRsWwtl
==
4'b0011
)
?
4'b0010
:
(
SVRsWwtl
==
4'b0100
)
?
4'b0110
:
(
SVRsWwtl
==
4'b0101
)
?
4'b0111
:
(
SVRsWwtl
==
4'b0110
)
?
4'b0101
:
(
SVRsWwtl
==
4'b0111
)
?
4'b0100
:
(
SVRsWwtl
==
4'b1000
)
?
4'b1100
:
(
SVRsWwtl
==
4'b1001
)
?
4'b1101
:
(
SVRsWwtl
==
4'b1010
)
?
4'b1111
:
(
SVRsWwtl
==
4'b1011
)
?
4'b1110
:
(
SVRsWwtl
==
4'b1100
)
?
4'b1010
:
(
SVRsWwtl
==
4'b1101
)
?
4'b1011
:
(
SVRsWwtl
==
4'b1110
)
?
4'b1001
:
4'b1000
;
reg
[
3
:
0
]
SVRomsOl
;
always
@
(
posedge
SVRHncAS
)
SVRomsOl
<=
SVReMSRP
;
initial
SVRomsOl
=
4'd0
;
reg
[
3
:
0
]
SVRtZEMw
,
SVRJzptl
;
always
@
(
posedge
SVRaNsOW
or
negedge
reset_n
)
if
(
~reset_n
)
SVRtZEMw
<=
4'd0
;
else
SVRtZEMw
<=
SVRomsOl
;
always
@
(
posedge
SVRaNsOW
or
negedge
reset_n
)
if
(
~reset_n
)
SVRJzptl
<=
4'd0
;
else
SVRJzptl
<=
SVRtZEMw
;
wire
[
3
:
0
]
SVRdGdCW
=
(
SVRJzptl
==
4'b0000
)
?
4'b0000
:
(
SVRJzptl
==
4'b0001
)
?
4'b0001
:
(
SVRJzptl
==
4'b0011
)
?
4'b0010
:
(
SVRJzptl
==
4'b0010
)
?
4'b0011
:
(
SVRJzptl
==
4'b0110
)
?
4'b0100
:
(
SVRJzptl
==
4'b0111
)
?
4'b0101
:
(
SVRJzptl
==
4'b0101
)
?
4'b0110
:
(
SVRJzptl
==
4'b0100
)
?
4'b0111
:
(
SVRJzptl
==
4'b1100
)
?
4'b1000
:
(
SVRJzptl
==
4'b1101
)
?
4'b1001
:
(
SVRJzptl
==
4'b1111
)
?
4'b1010
:
(
SVRJzptl
==
4'b1110
)
?
4'b1011
:
(
SVRJzptl
==
4'b1010
)
?
4'b1100
:
(
SVRJzptl
==
4'b1011
)
?
4'b1101
:
(
SVRJzptl
==
4'b1001
)
?
4'b1110
:
4'b1111
;
assign
SVRRgiPc
=
(
(
SVRjyLJF
^
SVRdGdCW
)
==
4'b0000
)
?
1'b1
:
1'b0
;
endmodule
module SVRzYBgZ
(
fclk
,
SVRJROZz
,
SVRcstsC
,
SVRfiOaI
,
SVRWNemH
,
SVRknyyH
,
SVRRZHEh
,
SVRySJvq
,
SVRpEcIs
,
SVRgAzyx
,
SVRcogji
,
SVRGGNIH
,
SVRhTMHu
,
SVRnaZWU
,
SVRfeSui
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRcstsC
;
input
SVRfiOaI
;
input
SVRWNemH
;
input
SVRknyyH
;
input
[
7
:
0
]
SVRRZHEh
;
input
SVRySJvq
;
input
[
5
:
0
]
SVRpEcIs
;
output
SVRgAzyx
;
output
SVRcogji
;
output
SVRGGNIH
;
output
SVRhTMHu
;
output
SVRnaZWU
;
output
SVRfeSui
;
wire
[
1
:
0
]
SVRnJxgP
;
assign
SVRnJxgP
=
{
SVRWNemH
,
SVRknyyH
}
;
parameter
SVRGRlDu
=
4'h0
;
parameter
SVRcPbhb
=
4'h1
;
parameter
SVRBUADa
=
4'h2
;
parameter
SVRzqjhR
=
4'h3
;
parameter
SVRmIEDV
=
4'h5
;
parameter
SVRgrPOX
=
4'h6
;
parameter
SVRPBQMp
=
4'h7
;
parameter
SVRghRLy
=
4'h8
;
parameter
SVRDDVsm
=
4'h9
;
parameter
SVRaITbX
=
4'hB
;
parameter
SVRmKstP
=
4'hC
;
parameter
SVRslfCl
=
4'hE
;
reg
[
7
:
0
]
SVRVyyGw
;
wire
[
7
:
0
]
SVRxmmqL
;
wire
SVRxZBAj
=
(
SVRVyyGw
>
SVRxmmqL
)
?
1'b1
:
1'b0
;
reg
[
3
:
0
]
SVRXSJFV
;
reg
[
3
:
0
]
SVRKPnIo
;
wire
SVReOCjy
;
wire
SVRcuOeM
;
wire
SVRbkuct
;
wire
SVRafkBJ
;
always
@
(
*
)
if
(
SVRcstsC
)
SVRKPnIo
=
SVRcPbhb
;
else
case
(
SVRXSJFV
)
SVRGRlDu
:
SVRKPnIo
=
SVRcPbhb
;
SVRcPbhb
:
if
(
(
SVRnJxgP
==
2'b11
)
&
SVRfiOaI
)
SVRKPnIo
=
SVRBUADa
;
else
SVRKPnIo
=
SVRcPbhb
;
SVRBUADa
:
if
(
SVRnJxgP
==
2'b01    // April-9-2015 manual change
)
SVRKPnIo
=
SVRzqjhR
;
else
SVRKPnIo
=
SVRBUADa
;
SVRzqjhR
:
if
(
SVRnJxgP
==
2'b00
)
SVRKPnIo
=
SVRmIEDV
;
else
if
(
SVRnJxgP
==
2'b11
)
SVRKPnIo
=
SVRBUADa
;
else
SVRKPnIo
=
SVRzqjhR
;
SVRmIEDV
:
begin
if
(
SVRxZBAj
==
1'b1
)
SVRKPnIo
=
SVRgrPOX
;
else
SVRKPnIo
=
SVRmIEDV
;
end
SVRgrPOX
:
begin
if
(
SVRxZBAj
==
1'b1
)
SVRKPnIo
=
SVRPBQMp
;
else
SVRKPnIo
=
SVRgrPOX
;
end
SVRPBQMp
:
begin
if
(
SVRySJvq
)
SVRKPnIo
=
SVRghRLy
;
else
SVRKPnIo
=
SVRPBQMp
;
end
SVRghRLy
:
begin
if
(
SVRnJxgP
!=
2'b00
)
SVRKPnIo
=
SVRDDVsm
;
else
SVRKPnIo
=
SVRghRLy
;
end
SVRDDVsm
:
begin
if
(
SVRnJxgP
==
2'b11
)
SVRKPnIo
=
SVRBUADa
;
else
if
(
SVRnJxgP
==
2'b00
)
SVRKPnIo
=
SVRghRLy
;
else
SVRKPnIo
=
SVRDDVsm
;
end
SVRaITbX
:
if
(
SVRnJxgP
==
2'b10
)
SVRKPnIo
=
SVRaITbX
;
else
if
(
SVRnJxgP
==
2'b00
)
SVRKPnIo
=
SVRmKstP
;
else
SVRKPnIo
=
SVRGRlDu
;
SVRmKstP
:
if
(
SVReOCjy
==
1'b1
)
SVRKPnIo
=
SVRslfCl
;
else
if
(
SVRbkuct
==
1'b1
)
SVRKPnIo
=
SVRGRlDu
;
else
if
(
SVRcuOeM
==
1'b1
)
SVRKPnIo
=
SVRGRlDu
;
else
SVRKPnIo
=
SVRmKstP
;
SVRslfCl
:
if
(
SVRnJxgP
==
2'b00
)
SVRKPnIo
=
SVRslfCl
;
else
SVRKPnIo
=
SVRGRlDu
;
default
:
SVRKPnIo
=
SVRGRlDu
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRXSJFV
<=
SVRGRlDu
;
else
if
(
SVRcstsC
==
1'b1
)
SVRXSJFV
<=
SVRcPbhb
;
else
SVRXSJFV
<=
SVRKPnIo
;
assign
SVRafkBJ
=
(
(
SVRXSJFV
==
SVRaITbX
)
&&
(
SVRKPnIo
==
SVRmKstP
)
)
?
1'b1
:
1'b0
;
SVRAcFNr
SVRnBPTi
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRcstsC
(
SVRcstsC
)
,
.SVRGNUwe
(
SVRnJxgP
[
1
]
)
,
.SVRcnTdT
(
SVRnJxgP
[
0
]
)
,
.SVRBGWBw
(
SVRafkBJ
)
,
.SVReOCjy
(
SVReOCjy
)
,
.SVRcuOeM
(
SVRcuOeM
)
,
.SVRbkuct
(
SVRbkuct
)
)
;
assign
SVRxmmqL
=
(
SVRXSJFV
==
SVRmIEDV
)
?
SVRRZHEh
:
(
SVRXSJFV
==
SVRgrPOX
)
?
{
2'h0
,
SVRpEcIs
}
:
8'h00
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRVyyGw
<=
8'h00
;
else
if
(
SVRcstsC
==
1'b1
)
SVRVyyGw
<=
8'h00
;
else
if
(
(
SVRXSJFV
==
SVRmIEDV
)
&
SVRxZBAj
)
SVRVyyGw
<=
8'h00
;
else
if
(
(
SVRXSJFV
!=
SVRmIEDV
)
&
(
SVRXSJFV
!=
SVRgrPOX
)
)
SVRVyyGw
<=
8'h00
;
else
SVRVyyGw
<=
SVRVyyGw
+
8'h01
;
reg
SVRcogji
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRcogji
<=
1'b0
;
else
if
(
SVRcstsC
==
1'b1
)
SVRcogji
<=
1'b0
;
else
if
(
SVRXSJFV
==
SVRPBQMp
)
SVRcogji
<=
1'b1
;
else
SVRcogji
<=
1'b0
;
assign
SVRgAzyx
=
(
SVRXSJFV
==
SVRghRLy
)
|
(
SVRKPnIo
==
SVRghRLy
)
|
(
SVRXSJFV
==
SVRDDVsm
)
;
assign
SVRGGNIH
=
(
SVRXSJFV
==
SVRPBQMp
)
|
(
SVRXSJFV
==
SVRghRLy
)
|
(
SVRXSJFV
==
SVRDDVsm
)
;
reg
SVRhTMHu
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRhTMHu
<=
1'b0
;
else
if
(
SVRXSJFV
==
SVRBUADa
)
SVRhTMHu
<=
1'b1
;
else
SVRhTMHu
<=
1'b0
;
reg
SVRnaZWU
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRnaZWU
<=
1'b0
;
else
if
(
SVRcstsC
==
1'b1
)
SVRnaZWU
<=
1'b0
;
else
if
(
(
SVRXSJFV
==
SVRghRLy
)
||
(
SVRXSJFV
==
SVRPBQMp
)
)
SVRnaZWU
<=
1'b1
;
else
SVRnaZWU
<=
1'b0
;
reg
SVRfeSui
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRfeSui
<=
1'b0
;
else
if
(
SVRcstsC
==
1'b1
)
SVRfeSui
<=
1'b0
;
else
if
(
SVRXSJFV
==
SVRGRlDu
)
SVRfeSui
<=
1'b1
;
else
SVRfeSui
<=
1'b0
;
endmodule
module SVRAcFNr
(
fclk
,
SVRJROZz
,
SVRcstsC
,
SVRGNUwe
,
SVRcnTdT
,
SVRBGWBw
,
SVReOCjy
,
SVRcuOeM
,
SVRbkuct
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRcstsC
;
input
SVRGNUwe
;
input
SVRcnTdT
;
input
SVRBGWBw
;
output
wire
SVReOCjy
;
output
wire
SVRcuOeM
;
output
wire
SVRbkuct
;
parameter
SVRnqYnL
=
8'h1e
;
parameter
SVRgiZGs
=
3'b000
;
parameter
SVRdEzqj
=
3'b100
;
parameter
SVRbPmIe
=
3'b101
;
parameter
SVRMnCjT
=
3'b110
;
parameter
SVRfakxn
=
3'b111
;
wire
[
1
:
0
]
SVRnJxgP
=
{
SVRGNUwe
,
SVRcnTdT
}
;
reg
[
2
:
0
]
SVRVoBcb
,
SVRoTaEX
;
always
@
(
SVRnJxgP
or
SVRBGWBw
or
SVRJROZz
or
SVReOCjy
or
SVRbkuct
or
SVRcuOeM
or
SVRVoBcb
)
case
(
SVRVoBcb
)
SVRgiZGs
:
if
(
SVRBGWBw
==
1'b1
)
SVRoTaEX
=
SVRdEzqj
;
else
SVRoTaEX
=
SVRgiZGs
;
SVRdEzqj
:
if
(
SVRBGWBw
==
1'b1
)
SVRoTaEX
=
SVRfakxn
;
else
if
(
SVRnJxgP
==
2'b10
)
SVRoTaEX
=
SVRMnCjT
;
else
if
(
SVRnJxgP
==
2'b01
)
SVRoTaEX
=
SVRbPmIe
;
else
if
(
SVRnJxgP
==
2'b00
)
SVRoTaEX
=
SVRdEzqj
;
else
SVRoTaEX
=
SVRfakxn
;
SVRbPmIe
:
if
(
SVRBGWBw
==
1'b1
)
SVRoTaEX
=
SVRfakxn
;
else
if
(
SVRnJxgP
==
2'b01
)
SVRoTaEX
=
SVRbPmIe
;
else
if
(
SVRnJxgP
==
2'b00
)
SVRoTaEX
=
SVRdEzqj
;
else
SVRoTaEX
=
SVRfakxn
;
SVRMnCjT
:
if
(
SVRBGWBw
==
1'b1
)
SVRoTaEX
=
SVRfakxn
;
else
if
(
SVRnJxgP
==
2'b10
)
SVRoTaEX
=
SVRMnCjT
;
else
if
(
SVRnJxgP
==
2'b00
)
SVRoTaEX
=
SVRdEzqj
;
else
SVRoTaEX
=
SVRfakxn
;
SVRfakxn
:
SVRoTaEX
=
SVRfakxn
;
default
:
SVRoTaEX
=
SVRfakxn
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRVoBcb
<=
SVRgiZGs
;
else
if
(
SVRcstsC
==
1'b1
)
SVRVoBcb
<=
SVRgiZGs
;
else
if
(
(
SVReOCjy
==
1'b1
)
||
(
SVRbkuct
==
1'b1
)
||
(
SVRcuOeM
==
1'b1
)
)
SVRVoBcb
<=
SVRgiZGs
;
else
SVRVoBcb
<=
SVRoTaEX
;
reg
[
3
:
0
]
SVRHwaPy
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRHwaPy
<=
4'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRcstsC
==
1'b1
)
===
1'bx
)
SVRHwaPy
<=
4'bxxxx
;
`endif
else
if
(
SVRcstsC
==
1'b1
)
SVRHwaPy
<=
4'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRoTaEX
==
SVRdEzqj
)
&&
(
(
SVRVoBcb
==
SVRbPmIe
)
||
(
SVRVoBcb
==
SVRMnCjT
)
)
)
===
1'bx
)
SVRHwaPy
<=
4'bxxxx
;
`endif
else
if
(
(
SVRoTaEX
==
SVRdEzqj
)
&&
(
(
SVRVoBcb
==
SVRbPmIe
)
||
(
SVRVoBcb
==
SVRMnCjT
)
)
)
SVRHwaPy
<=
SVRHwaPy
+
4'd1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVReOCjy
==
1'b1
)
||
(
SVRbkuct
==
1'b1
)
||
(
SVRcuOeM
==
1'b1
)
)
===
1'bx
)
SVRHwaPy
<=
4'bxxx
;
`endif
else
if
(
(
SVReOCjy
==
1'b1
)
||
(
SVRbkuct
==
1'b1
)
||
(
SVRcuOeM
==
1'b1
)
)
SVRHwaPy
<=
3'd0
;
reg
[
7
:
0
]
SVRqlAum
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRqlAum
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRcstsC
==
1'b1
)
===
1'bx
)
SVRqlAum
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRcstsC
==
1'b1
)
SVRqlAum
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRHwaPy
==
4'd9
)
===
1'bx
)
SVRqlAum
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRHwaPy
==
4'd9
)
SVRqlAum
<=
SVRqlAum
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRoTaEX
==
SVRMnCjT
)
&&
(
SVRVoBcb
==
SVRdEzqj
)
)
===
1'bx
)
SVRqlAum
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRoTaEX
==
SVRMnCjT
)
&&
(
SVRVoBcb
==
SVRdEzqj
)
)
SVRqlAum
<=
{
SVRqlAum
[
6
:
0
]
,
1'b1
}
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRoTaEX
==
SVRbPmIe
)
&&
(
SVRVoBcb
==
SVRdEzqj
)
)
===
1'bx
)
SVRqlAum
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRoTaEX
==
SVRbPmIe
)
&&
(
SVRVoBcb
==
SVRdEzqj
)
)
SVRqlAum
<=
{
SVRqlAum
[
6
:
0
]
,
1'b0
}
;
assign
SVReOCjy
=
(
SVRHwaPy
!=
4'd9
)
?
1'b0
:
(
SVRVoBcb
==
SVRfakxn
)
?
1'b0
:
(
SVRqlAum
==
SVRnqYnL
)
?
1'b1
:
1'b0
;
assign
SVRbkuct
=
(
SVRHwaPy
!=
4'd9
)
?
1'b0
:
(
SVRVoBcb
==
SVRfakxn
)
?
1'b0
:
(
SVRqlAum
==
SVRnqYnL
)
?
1'b0
:
1'b1
;
assign
SVRcuOeM
=
(
SVRVoBcb
==
SVRfakxn
)
?
1'b1
:
1'b0
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRuPrNG
(
fclk
,
SVRJROZz
,
SVRcstsC
,
SVRfiOaI
,
SVRWNemH
,
SVRknyyH
,
SVRRZHEh
,
SVRGGNIH
,
SVRhTMHu
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRcstsC
;
input
SVRfiOaI
;
input
SVRWNemH
;
input
SVRknyyH
;
input
[
7
:
0
]
SVRRZHEh
;
output
SVRGGNIH
;
output
SVRhTMHu
;
reg
[
7
:
0
]
SVRVyyGw
;
wire
SVRxZBAj
;
wire
[
1
:
0
]
SVRnJxgP
;
assign
SVRnJxgP
=
{
SVRWNemH
,
SVRknyyH
}
;
parameter
SVRBUADa
=
2'd0
;
parameter
SVRsdNEU
=
2'd2
;
parameter
SVRghRLy
=
2'd3
;
reg
[
1
:
0
]
SVRKPnIo
;
reg
[
1
:
0
]
SVRXSJFV
;
always
@
(
*
)
case
(
SVRXSJFV
)
SVRBUADa
:
if
(
SVRnJxgP
==
2'b00
)
SVRKPnIo
=
SVRsdNEU
;
else
SVRKPnIo
=
SVRBUADa
;
SVRsdNEU
:
if
(
SVRxZBAj
==
1'b1
)
SVRKPnIo
=
SVRghRLy
;
else
SVRKPnIo
=
SVRsdNEU
;
SVRghRLy
:
if
(
SVRnJxgP
!=
2'b00
)
SVRKPnIo
=
SVRBUADa
;
else
SVRKPnIo
=
SVRghRLy
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRXSJFV
<=
SVRBUADa
;
else
if
(
SVRcstsC
==
1'b1
)
SVRXSJFV
<=
SVRBUADa
;
else
SVRXSJFV
<=
SVRKPnIo
;
assign
SVRxZBAj
=
(
SVRVyyGw
>=
SVRRZHEh
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRVyyGw
<=
8'h00
;
else
if
(
SVRcstsC
==
1'b1
)
SVRVyyGw
<=
8'h00
;
else
if
(
(
SVRXSJFV
!=
SVRsdNEU
)
)
SVRVyyGw
<=
8'h00
;
else
SVRVyyGw
<=
SVRVyyGw
+
8'h01
;
assign
SVRGGNIH
=
(
SVRXSJFV
==
SVRghRLy
)
;
wire
SVRhTMHu
=
(
SVRXSJFV
==
SVRBUADa
)
?
1'b1
:
1'b0
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRDWPuG
(
SVRcstsC
,
SVRfSoOm
,
fclk
,
pclk
,
SVRrGCzn
,
SVRzMTVm
,
SVRWiNOI
,
SVRyEtuR
,
SVRyMsqX
,
SVRmtjIy
,
SVRSCAjD
,
SVRhzkfv
,
SVRuPKrP
,
SVRYgHNS
,
SVRWnoBL
,
SVRLwmmN
,
SVRVYyIN
,
SVRJsIJK
,
SVRopDmx
,
SVROEvJE
,
SVRnCFbF
,
svr_pixel
,
svr_pixel_valid
,
SVRgDTYn
,
svr_fs
,
svr_fe
,
svr_ls
,
svr_le
,
svr_data_type
,
svr_cpu_int
,
SVRTVbtZ
,
SVRHXUZw
,
SVRZyNzG
,
SVRCqyoW
,
SVRDmFCK
,
SVRjFeTQ
,
SVRIgOeF
,
SVRQiYom
,
SVRTAKyC
,
SVRUxrba
)
;
input
SVRcstsC
;
output
SVRfSoOm
;
input
fclk
;
input
pclk
;
input
SVRrGCzn
;
input
SVRzMTVm
;
input
SVRWiNOI
;
input
SVRyEtuR
;
input
[
5
:
0
]
SVRyMsqX
;
input
[
31
:
0
]
SVRmtjIy
;
input
SVRSCAjD
;
input
[
7
:
0
]
SVRhzkfv
;
input
SVRuPKrP
;
input
SVRYgHNS
;
input
SVRWnoBL
;
input
SVRLwmmN
;
input
SVRVYyIN
;
input
SVRJsIJK
;
input
SVRopDmx
;
input
SVROEvJE
;
input
SVRnCFbF
;
output
[
23
:
0
]
svr_pixel
;
output
svr_pixel_valid
;
output
[
1
:
0
]
SVRgDTYn
;
output
svr_fs
;
output
svr_fe
;
output
svr_ls
;
output
svr_le
;
`ifdef SVRyllEh 
output
SVRMFfPD
;
output
SVRTPCUO
;
`endif
output
[
5
:
0
]
svr_data_type
;
output
svr_cpu_int
;
output
[
31
:
0
]
SVRTVbtZ
;
output
[
27
:
0
]
SVRHXUZw
;
output
SVRZyNzG
;
`ifdef SVRsQYvh 
output
[
31
:
0
]
SVRioKpl
;
`endif
`ifdef SVRCadQw 
output
SVRCqyoW
;
input
[
7
:
0
]
SVRDmFCK
;
input
SVRjFeTQ
;
input
SVRIgOeF
;
input
SVRQiYom
;
input
SVRTAKyC
;
input
SVRUxrba
;
`endif
wire
SVRehSHF
;
wire
[
31
:
0
]
SVRCdWQP
;
wire
[
5
:
0
]
SVRaVTNl
;
wire
SVRMQsMw
;
wire
SVRFoFlc
;
wire
SVRBAlYr
;
wire
SVRzGBRz
;
wire
SVRmQNVM
;
wire
SVRgVTxt
;
wire
[
31
:
0
]
SVRDXWLJ
;
wire
[
31
:
0
]
SVRasuLi
;
wire
[
31
:
0
]
SVRmcglv
;
assign
SVRzGBRz
=
1'b1
;
assign
SVRmQNVM
=
1'b0
;
assign
SVRgVTxt
=
1'b0
;
wire
SVRZyNzG
=
SVRMQsMw
&
SVRzGBRz
;
SVRgbDFk
SVRPtkiW
(
.fclk
(
fclk
)
,
.pclk
(
pclk
)
,
.SVRJROZz
(
SVRWiNOI
)
,
.SVRgdBWO
(
SVRrGCzn
)
,
.SVRDBnyu
(
SVRzMTVm
)
,
.SVRmtjIy
(
SVRmtjIy
)
,
.SVRCdWQP
(
SVRCdWQP
)
,
.address
(
SVRyMsqX
)
,
.SVRaVTNl
(
SVRaVTNl
)
,
.SVRSCAjD
(
SVRSCAjD
)
,
.SVRehSHF
(
SVRehSHF
)
)
;
wire
[
27
:
0
]
SVRUtdgF
;
wire
[
27
:
0
]
SVRHXUZw
;
wire
[
31
:
0
]
SVRjDxvg
;
assign
SVRjDxvg
[
14
]
=
1'b0
;
assign
SVRjDxvg
[
13
]
=
1'b0
;
assign
SVRjDxvg
[
12
]
=
1'b0
;
assign
SVRjDxvg
[
11
]
=
1'b0
;
assign
SVRjDxvg
[
10
]
=
1'b1
;
assign
SVRjDxvg
[
9
]
=
1'b0
;
assign
SVRjDxvg
[
8
]
=
1'b0
;
assign
SVRjDxvg
[
7
]
=
SVRQiYom
;
assign
SVRjDxvg
[
6
]
=
SVRJsIJK
;
assign
SVRjDxvg
[
5
]
=
SVRVYyIN
;
assign
SVRjDxvg
[
6
]
=
SVRJsIJK
;
assign
SVRjDxvg
[
4
]
=
1'b0
;
assign
SVRjDxvg
[
3
]
=
1'b0
;
assign
SVRjDxvg
[
2
]
=
SVRIgOeF
;
assign
SVRjDxvg
[
1
]
=
SVRYgHNS
;
assign
SVRjDxvg
[
0
]
=
SVRWnoBL
;
wire
[
1
:
0
]
SVREOLkD
;
wire
[
31
:
0
]
SVRBNOxF
;
wire
[
31
:
0
]
SVRZmqEG
;
wire
[
15
:
0
]
SVRLZDhh
;
wire
[
15
:
0
]
SVReTkwu
;
wire
[
15
:
0
]
SVROpBdB
;
wire
SVRUHNBN
;
wire
SVRXQTNt
;
wire
SVRyVWTJ
;
wire
SVRMxYWr
;
wire
SVRTlzYi
;
wire
[
7
:
0
]
SVRWFmze
;
wire
[
7
:
0
]
SVRkjcfT
;
wire
SVRRXWun
;
wire
SVRVyyKg
;
wire
[
15
:
0
]
SVRxmmsd
;
wire
[
7
:
0
]
SVRxZBBs
;
wire
[
31
:
0
]
SVRXSjgA
;
wire
SVRKPAVd
;
wire
SVReojQs
;
wire
SVRoAAnA
;
wire
SVRhnNgN
;
wire
SVRDGtDt
;
wire
SVRoQJOJ
;
wire
[
15
:
0
]
SVRhVrUr
;
wire
SVRPQEPZ
;
wire
SVRGolNq
;
wire
SVRCAbmZ
;
wire
[
31
:
0
]
SVRoNaGz
;
wire
[
31
:
0
]
SVRTmwId
;
wire
[
31
:
0
]
SVRwglRb
;
wire
[
31
:
0
]
SVRxwbOR
;
wire
[
31
:
0
]
SVRlLaUV
;
wire
[
31
:
0
]
SVRFsaXX
;
wire
SVRBcWQp
;
assign
SVRfSoOm
=
SVRUtdgF
[
0
]
;
wire
SVRLljSa
;
assign
SVRLljSa
=
SVRZyNzG
;
wire
SVRzUTNy
=
SVRcstsC
;
wire
[
23
:
0
]
SVRyQsmd
;
wire
SVRmvjGB
;
wire
[
5
:
0
]
SVRGKeQn
;
wire
[
23
:
0
]
SVRqscVG
;
wire
SVRucXph
;
assign
svr_pixel
=
(
SVRmQNVM
)
?
SVRyQsmd
:
SVRqscVG
;
assign
svr_pixel_valid
=
(
SVRmQNVM
)
?
SVRmvjGB
:
SVRucXph
;
SVRwuuAu
SVRlkknk
(
.SVRJROZz
(
SVRyEtuR
)
,
.fclk
(
fclk
)
,
.SVRrYaZV
(
SVRyQsmd
[
23
:
0
]
)
,
.SVRizAZX
(
SVRmvjGB
)
,
.SVRQfjSP
(
svr_ls
)
,
.SVRhwAOL
(
svr_fs
)
,
.SVRdlnUs
(
SVRqscVG
[
23
:
0
]
)
,
.SVRBFgxj
(
SVRucXph
)
)
;
reg
[
1
:
0
]
SVRLxvHB
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRLxvHB
<=
2'b00
;
else
SVRLxvHB
<=
SVRUtdgF
[
2
:
1
]
;
`ifdef SVRCadQw 
assign
SVRCqyoW
=
(
SVRLxvHB
==
2'b00
)
?
1'b0
:
1'b1
;
`endif
`ifdef SVReFgJe 
assign
SVRCpDrC
=
SVRLxvHB
[
1
]
;
`endif
`ifdef SVRaBkbf 
assign
SVRMgbtT
=
(
SVRLxvHB
==
2'b11
)
?
1'b1
:
1'b0
;
`endif
SVRFwWBn
SVRBeuGx
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRLwmmN
(
SVRLwmmN
)
,
.SVRnckQL
(
SVRLZDhh
[
15
:
0
]
)
,
.SVRsUANj
(
SVRXQTNt
)
,
.SVRhzkfv
(
SVRhzkfv
[
7
:
0
]
)
,
.SVRuPKrP
(
SVRuPKrP
)
,
.SVRJsIJK
(
SVRJsIJK
)
,
.SVRvqjMV
(
SVRRXWun
)
`ifdef SVRCadQw 
,
.SVRCqyoW
(
SVRCqyoW
)
,
.SVRDmFCK
(
SVRDmFCK
[
7
:
0
]
)
,
.SVRjFeTQ
(
SVRjFeTQ
)
,
.SVRQiYom
(
SVRQiYom
)
`endif
`ifdef SVReFgJe 
,
.SVRCpDrC
(
SVRCpDrC
)
,
.SVRwBALo
(
SVRwBALo
[
7
:
0
]
)
,
.SVRLnNsH
(
SVRLnNsH
)
,
.SVRSGtJq
(
SVRSGtJq
)
`endif
`ifdef SVRaBkbf 
,
.SVRMgbtT
(
SVRMgbtT
)
,
.SVRIJfkz
(
SVRIJfkz
[
7
:
0
]
)
,
.SVRdLyxD
(
SVRdLyxD
)
,
.SVRNliEf
(
SVRNliEf
)
`endif
)
;
SVRfZzHt
SVROSiJA
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRGpakE
(
SVRLZDhh
[
15
:
0
]
)
,
.SVRcbwXF
(
SVRXQTNt
)
,
.SVRBaLYP
(
SVReTkwu
[
15
:
0
]
)
,
.SVRnAsZu
(
SVRyVWTJ
)
,
.SVRMxYWr
(
SVRMxYWr
)
,
.SVRsgfsB
(
SVRRXWun
)
,
.SVRvwyBE
(
SVRUtdgF
[
4
]
)
,
.SVRPQEPZ
(
SVRPQEPZ
)
,
.SVRGolNq
(
SVRGolNq
)
,
.SVRCAbmZ
(
SVRCAbmZ
)
,
.SVRhVrUr
(
SVRhVrUr
[
15
:
0
]
)
,
.SVRklMnp
(
SVRWFmze
[
7
:
0
]
)
,
.SVRFfTGh
(
SVRTlzYi
)
,
.SVRbwSIu
(
SVRKPAVd
)
)
;
SVRalwrK
SVRMYgbJ
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRFoFlc
(
SVRFoFlc
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVRyMsqX
(
SVRaVTNl
)
,
.SVRmtjIy
(
SVRCdWQP
[
31
:
0
]
)
,
.SVRUtdgF
(
SVRUtdgF
[
16
:
5
]
)
,
.SVRGolNq
(
SVRGolNq
)
,
.SVRCAbmZ
(
SVRCAbmZ
)
,
.SVRhVrUr
(
SVRhVrUr
[
15
:
0
]
)
,
.SVRFsZsI
(
SVRWFmze
[
7
:
0
]
)
,
.SVRBCVbi
(
SVRKPAVd
)
,
.SVRnOXaE
(
SVReTkwu
[
15
:
0
]
)
,
.SVRcbwXF
(
SVRyVWTJ
)
,
.SVRMxYWr
(
SVRMxYWr
)
,
.SVRBaLYP
(
SVROpBdB
[
15
:
0
]
)
,
.SVRnAsZu
(
SVRUHNBN
)
,
.SVRBcWQp
(
SVRBcWQp
)
,
.SVRgUyap
(
SVRkjcfT
[
7
:
0
]
)
,
.SVRpqIsy
(
SVReojQs
)
,
.SVRsgfsB
(
SVRTlzYi
)
,
.SVRhirjM
(
SVRVyyKg
)
,
.SVRvwyBE
(
SVRUtdgF
[
4
]
)
,
.SVRpxeXJ
(
SVRjDxvg
[
1
]
)
,
.SVRHlCYR
(
SVRjDxvg
[
30
]
)
,
.SVRQfoZV
(
SVRjDxvg
[
29
]
)
,
.SVREOLkD
(
SVREOLkD
[
1
:
0
]
)
,
.SVRBNOxF
(
SVRBNOxF
[
31
:
0
]
)
,
.SVRhWcSo
(
SVRoAAnA
)
,
.SVRxmmsd
(
SVRxmmsd
[
15
:
0
]
)
,
.SVRDGtDt
(
SVRDGtDt
)
,
.SVRhnNgN
(
SVRhnNgN
)
,
.SVRGKeQn
(
SVRGKeQn
)
,
.SVRBAlYr
(
SVRBAlYr
)
)
;
`ifdef SVRprxoy 
SVRTBHZc
SVRWNQzB
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRknrFe
(
SVROpBdB
[
15
:
0
]
)
,
.SVRsUANj
(
SVRUHNBN
)
,
.SVRRzeiT
(
SVRkjcfT
[
5
:
0
]
)
,
.SVRoAAnA
(
SVRoAAnA
)
,
.SVRVmcEw
(
SVRyQsmd
[
23
:
0
]
)
,
.SVRGKeQn
(
SVRGKeQn
)
,
.SVRUtdgF
(
SVRUtdgF
[
27
:
0
]
)
,
.SVRxgbpl
(
SVRmvjGB
)
,
.SVRoQJOJ
(
SVRoQJOJ
)
,
.SVRBcWQp
(
SVRBcWQp
)
,
.SVRlDAHF
(
svr_ls
)
)
;
`endif
`ifndef SVRprxoy
SVRFoNQp
SVRWNQzB
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRknrFe
(
SVROpBdB
[
15
:
0
]
)
,
.SVRsUANj
(
SVRUHNBN
)
,
.SVRBcWQp
(
SVRBcWQp
)
,
.SVRoAAnA
(
SVRoAAnA
)
,
.SVRVmcEw
(
SVRyQsmd
[
23
:
0
]
)
,
.SVRGKeQn
(
SVRGKeQn
)
,
.SVRxgbpl
(
SVRmvjGB
)
,
.SVRoQJOJ
(
SVRoQJOJ
)
)
;
`endif
SVRBAPNY
SVRzGqmq
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRFoFlc
(
SVRFoFlc
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVRyMsqX
(
SVRaVTNl
)
,
.SVRmtjIy
(
SVRCdWQP
[
28
:
15
]
)
,
.SVRmqigi
(
SVRUtdgF
[
0
]
)
,
.SVRLljSa
(
SVRLljSa
)
,
.SVRYgHNS
(
SVRYgHNS
)
,
.SVRopDmx
(
SVRopDmx
)
,
.SVROEvJE
(
SVROEvJE
)
,
.SVRCqyoW
(
SVRCqyoW
)
,
.SVRTAKyC
(
SVRTAKyC
)
,
.SVRUxrba
(
SVRUxrba
)
,
.SVRnCFbF
(
SVRnCFbF
)
,
.SVRjDxvg
(
SVRjDxvg
[
31
:
15
]
)
)
;
SVRsbAVU
SVRJaNxX
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRFoFlc
(
SVRFoFlc
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVRyMsqX
(
SVRaVTNl
)
,
.SVRDtpEP
(
SVRCdWQP
[
31
:
17
]
)
,
.SVROJhPU
(
SVRCdWQP
[
7
:
0
]
)
,
.SVREOLkD
(
SVREOLkD
[
1
:
0
]
)
,
.SVRBNOxF
(
SVRBNOxF
[
30
:
29
]
)
,
.SVRklMnp
(
SVRkjcfT
[
7
:
0
]
)
,
.SVRbwSIu
(
SVReojQs
)
,
.SVRvwyBE
(
SVRUtdgF
[
4
]
)
,
.SVRPQEPZ
(
SVRPQEPZ
)
,
.SVRGolNq
(
SVRGolNq
)
,
.SVRCAbmZ
(
SVRCAbmZ
)
,
.SVRZmqEG
(
SVRZmqEG
[
31
:
0
]
)
,
.SVRDGtDt
(
SVRDGtDt
)
,
.SVRhnNgN
(
SVRhnNgN
)
)
;
SVRURDuX
SVRjPKCp
(
.fclk
(
fclk
)
,
.pclk
(
pclk
)
,
.SVRyEtuR
(
SVRyEtuR
)
,
.SVRWiNOI
(
SVRWiNOI
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRrGCzn
(
SVRrGCzn
)
,
.SVRzMTVm
(
SVRzMTVm
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVREusOH
(
SVRaVTNl
)
,
.SVRBdFMH
(
SVRyMsqX
)
,
.SVRmtjIy
(
SVRCdWQP
[
31
:
0
]
)
,
.SVRSCAjD
(
SVRSCAjD
)
,
.SVRklMnp
(
SVRkjcfT
[
7
:
0
]
)
,
.SVRjDxvg
(
SVRjDxvg
[
30
:
29
]
)
,
.SVREOLkD
(
SVREOLkD
[
1
:
0
]
)
,
.SVRZmqEG
(
SVRZmqEG
[
30
:
28
]
)
,
.SVRBNOxF
(
SVRBNOxF
[
30
:
29
]
)
,
.SVRxmmsd
(
SVRxmmsd
[
15
:
0
]
)
,
.SVRbwSIu
(
SVReojQs
)
,
.SVRxZBBs
(
SVRxZBBs
[
7
:
0
]
)
,
.SVRXSjgA
(
SVRXSjgA
[
31
:
0
]
)
,
.SVRFoFlc
(
SVRFoFlc
)
,
.svr_cpu_int
(
svr_cpu_int
)
)
;
SVRZuLLH
SVRLDoLh
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVRyMsqX
(
SVRaVTNl
)
,
.SVRmtjIy
(
SVRCdWQP
)
,
.SVRUtdgF
(
SVRUtdgF
[
27
:
0
]
)
,
.SVRHXUZw
(
SVRHXUZw
[
27
:
0
]
)
,
.SVRSoHSD
(
SVRDXWLJ
)
,
.SVRwHqWo
(
SVRasuLi
)
,
.SVRXjEqy
(
SVRmcglv
)
)
;
SVRkYKaD
SVRfzsAo
(
.fclk
(
fclk
)
,
.pclk
(
pclk
)
,
.SVRyEtuR
(
SVRyEtuR
)
,
.SVRWiNOI
(
SVRWiNOI
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRrGCzn
(
SVRrGCzn
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVREusOH
(
SVRaVTNl
)
,
.SVRBdFMH
(
SVRyMsqX
)
,
.SVRCmjnh
(
SVRCdWQP
[
0
]
)
,
.SVRSCAjD
(
SVRSCAjD
)
,
.SVRgVTxt
(
SVRgVTxt
)
,
.SVRUtdgF
(
SVRUtdgF
[
27
:
0
]
)
,
.SVRHXUZw
(
SVRHXUZw
[
27
:
0
]
)
,
.SVRxZBBs
(
SVRxZBBs
[
7
:
0
]
)
,
.SVRXSjgA
(
SVRXSjgA
[
31
:
0
]
)
,
.SVRjDxvg
(
SVRjDxvg
[
31
:
0
]
)
,
.SVREOLkD
(
SVREOLkD
[
1
:
0
]
)
,
.SVRBNOxF
(
SVRBNOxF
[
31
:
0
]
)
,
.SVRZmqEG
(
SVRZmqEG
[
31
:
0
]
)
,
.SVRoQJOJ
(
SVRoQJOJ
)
,
.SVRAzazu
(
SVRMxYWr
)
,
.SVRklMnp
(
SVRkjcfT
[
7
:
0
]
)
,
.SVRbwSIu
(
SVReojQs
)
,
.SVRZfWeB
(
SVRVyyKg
)
,
.SVRTVbtZ
(
SVRTVbtZ
[
31
:
0
]
)
,
.SVRZyNzG
(
SVRMQsMw
)
,
.SVRgDTYn
(
SVRgDTYn
)
,
.svr_fs
(
svr_fs
)
,
.svr_fe
(
svr_fe
)
,
.svr_ls
(
svr_ls
)
,
.svr_le
(
svr_le
)
,
`ifdef SVRyllEh 
.SVRMFfPD
(
SVRMFfPD
)
,
.SVRTPCUO
(
SVRTPCUO
)
,
`endif
.svr_data_type
(
svr_data_type
[
5
:
0
]
)
`ifdef SVRNJLgb 
,
.SVRoNaGz
(
SVRoNaGz
[
31
:
0
]
)
,
.SVRTmwId
(
SVRTmwId
[
31
:
0
]
)
,
.SVRwglRb
(
SVRwglRb
[
31
:
0
]
)
,
.SVRxwbOR
(
SVRxwbOR
[
31
:
0
]
)
,
.SVRlLaUV
(
SVRlLaUV
[
31
:
0
]
)
,
.SVRFsaXX
(
SVRFsaXX
[
31
:
0
]
)
`endif
)
;
`ifdef SVRNJLgb 
SVRlWTue
SVRfYwkC
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRyEtuR
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRehSHF
(
SVRehSHF
)
,
.SVRyMsqX
(
SVRaVTNl
)
,
.SVRmtjIy
(
SVRCdWQP
[
31
:
0
]
)
,
.SVRopDmx
(
SVRopDmx
)
,
.SVRTAKyC
(
SVRTAKyC
)
,
.SVRczlfo
(
SVRBAlYr
)
,
.SVRGolNq
(
SVRGolNq
)
,
.SVRCAbmZ
(
SVRCAbmZ
)
,
.SVRoNaGz
(
SVRoNaGz
[
31
:
0
]
)
,
.SVRTmwId
(
SVRTmwId
[
31
:
0
]
)
,
.SVRwglRb
(
SVRwglRb
[
31
:
0
]
)
,
.SVRxwbOR
(
SVRxwbOR
[
31
:
0
]
)
,
.SVRlLaUV
(
SVRlLaUV
[
31
:
0
]
)
,
.SVRFsaXX
(
SVRFsaXX
[
31
:
0
]
)
)
;
`endif
endmodule
module SVRgbDFk
(
fclk
,
pclk
,
SVRJROZz
,
SVRgdBWO
,
SVRDBnyu
,
SVRSCAjD
,
SVRmtjIy
,
address
,
SVRaVTNl
,
SVRCdWQP
,
SVRehSHF
)
;
input
fclk
;
input
pclk
;
input
SVRJROZz
;
input
SVRgdBWO
;
input
SVRDBnyu
;
input
SVRSCAjD
;
input
[
31
:
0
]
SVRmtjIy
;
input
[
5
:
0
]
address
;
output
[
5
:
0
]
SVRaVTNl
;
output
[
31
:
0
]
SVRCdWQP
;
output
SVRehSHF
;
reg
SVRRqewu
;
reg
[
31
:
0
]
SVRCdWQP
;
reg
[
5
:
0
]
SVRaVTNl
;
initial
#
0
SVRRqewu
=
1'b0
;
always
@
(
posedge
pclk
)
if
(
(
SVRDBnyu
==
1'b1
)
&&
(
SVRgdBWO
==
1'b1
)
&&
(
SVRSCAjD
==
1'b1
)
)
SVRRqewu
<=
1'b1
;
else
SVRRqewu
<=
1'b0
;
wire
SVRviclk
=
(
SVRDBnyu
&
SVRgdBWO
&
SVRSCAjD
&
(
~SVRRqewu
)
)
;
initial
#
0
SVRaVTNl
=
6'd0
;
always
@
(
posedge
pclk
)
if
(
SVRviclk
)
SVRaVTNl
<=
address
;
initial
#
0
SVRCdWQP
=
32'd0
;
always
@
(
posedge
pclk
)
if
(
SVRviclk
)
SVRCdWQP
<=
SVRmtjIy
;
wire
SVRwXWXv
;
reg
SVRXruRB
;
initial
#
0
SVRXruRB
=
1'b0
;
always
@
(
posedge
pclk
)
if
(
SVRwXWXv
)
SVRXruRB
<=
1'b0
;
else
if
(
SVRviclk
)
SVRXruRB
<=
1'b1
;
wire
SVRkcgOe
,
SVRfbduC
;
SVRRWXII
SVRCAbko
(
.SVRSrADr
(
SVRkcgOe
)
,
.SVRnXiwb
(
SVRXruRB
)
,
.SVRlqCbq
(
fclk
)
)
;
SVRRWXII
SVRoNafH
(
.SVRSrADr
(
SVRfbduC
)
,
.SVRnXiwb
(
SVRkcgOe
)
,
.SVRlqCbq
(
fclk
)
)
;
wire
SVRTmWuh
,
SVRwgyKD
;
SVRRWXII
SVRxWHKF
(
.SVRSrADr
(
SVRTmWuh
)
,
.SVRnXiwb
(
SVRfbduC
)
,
.SVRlqCbq
(
pclk
)
)
;
SVRRWXII
SVRxRMKG
(
.SVRSrADr
(
SVRwgyKD
)
,
.SVRnXiwb
(
SVRTmWuh
)
,
.SVRlqCbq
(
pclk
)
)
;
assign
SVRwXWXv
=
SVRwgyKD
;
reg
SVRXoPkh
;
initial
#
0
SVRXoPkh
=
1'b0
;
always
@
(
posedge
fclk
)
SVRXoPkh
<=
SVRfbduC
;
assign
SVRehSHF
=
(
(
~SVRXoPkh
)
&
SVRfbduC
)
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRlWTue
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRehSHF
,
SVRyMsqX
,
SVRmtjIy
,
SVRopDmx
,
SVRTAKyC
,
SVRczlfo
,
SVRGolNq
,
SVRCAbmZ
,
SVRoNaGz
,
SVRTmwId
,
SVRwglRb
,
SVRxwbOR
,
SVRlLaUV
,
SVRFsaXX
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRzUTNy
;
input
SVRehSHF
;
input
[
7
:
2
]
SVRyMsqX
;
input
[
31
:
0
]
SVRmtjIy
;
input
SVRopDmx
;
input
SVRTAKyC
;
input
SVRczlfo
;
input
SVRGolNq
;
input
SVRCAbmZ
;
output
[
31
:
0
]
SVRoNaGz
;
output
[
31
:
0
]
SVRTmwId
;
output
[
31
:
0
]
SVRwglRb
;
output
[
31
:
0
]
SVRxwbOR
;
output
[
31
:
0
]
SVRlLaUV
;
output
[
31
:
0
]
SVRFsaXX
;
reg
[
31
:
0
]
SVRVyyGw
;
reg
[
31
:
0
]
SVRfJLFv
;
reg
[
31
:
0
]
SVROKoIB
;
reg
[
31
:
0
]
SVRGlDJE
;
reg
[
31
:
0
]
SVRczkkG
;
reg
[
31
:
0
]
SVRBmffQ
;
reg
SVRnGCcv
;
reg
[
9
:
0
]
SVRgqoBK
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRgqoBK
<=
10'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRgqoBK
<=
10'bxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRgqoBK
<=
10'd0
;
else
SVRgqoBK
<=
SVRgqoBK
+
10'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRVyyGw
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRgnUJW
)
)
===
1'bx
)
SVRVyyGw
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRgnUJW
)
)
SVRVyyGw
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRVyyGw
!=
32'd0
)
&&
(
SVRgqoBK
==
10'h3ff
)
)
===
1'bx
)
SVRVyyGw
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRVyyGw
!=
32'd0
)
&&
(
SVRgqoBK
==
10'h3ff
)
&&
(
~SVRzUTNy
)
)
SVRVyyGw
<=
SVRVyyGw
+
32'hffffffff
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRnGCcv
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRnGCcv
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRnGCcv
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRVyyGw
!=
32'd0
)
===
1'bx
)
SVRnGCcv
<=
1'bx
;
`endif
else
if
(
SVRVyyGw
!=
32'd0
)
SVRnGCcv
<=
1'b1
;
else
SVRnGCcv
<=
1'b0
;
reg
SVRdiHns
;
reg
SVRnxmZZ
;
reg
SVRGlGZz
;
reg
SVRcZlSD
;
reg
SVRNSBOF
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRdiHns
<=
1'b0
;
else
SVRdiHns
<=
SVRopDmx
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRnxmZZ
<=
1'b0
;
else
SVRnxmZZ
<=
SVRTAKyC
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRGlGZz
<=
1'b0
;
else
SVRGlGZz
<=
SVRczlfo
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRcZlSD
<=
1'b0
;
else
SVRcZlSD
<=
SVRGolNq
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRNSBOF
<=
1'b0
;
else
SVRNSBOF
<=
SVRCAbmZ
;
reg
SVRFPJMg
;
reg
SVRbONlu
;
reg
SVRmNpYA
;
reg
SVRSMDrE
;
reg
SVRwTOiP
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRFPJMg
<=
1'b0
;
else
SVRFPJMg
<=
(
SVRopDmx
&
~
SVRdiHns
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRbONlu
<=
1'b0
;
else
SVRbONlu
<=
(
SVRTAKyC
&
~
SVRnxmZZ
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRmNpYA
<=
1'b0
;
else
SVRmNpYA
<=
(
SVRczlfo
&
~
SVRGlGZz
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRSMDrE
<=
1'b0
;
else
SVRSMDrE
<=
(
SVRGolNq
&
~
SVRcZlSD
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRwTOiP
<=
1'b0
;
else
SVRwTOiP
<=
(
SVRCAbmZ
&
~
SVRNSBOF
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRfJLFv
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRfJLFv
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRfJLFv
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRPZskp
)
)
===
1'bx
)
SVRfJLFv
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRPZskp
)
)
SVRfJLFv
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRFPJMg
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRfJLFv
!=
32'hffffffff
)
)
===
1'bx
)
SVRfJLFv
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRFPJMg
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRfJLFv
!=
32'hffffffff
)
)
SVRfJLFv
<=
SVRfJLFv
+
32'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVROKoIB
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVROKoIB
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVROKoIB
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRgtFxy
)
)
===
1'bx
)
SVROKoIB
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRgtFxy
)
)
SVROKoIB
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRbONlu
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVROKoIB
!=
32'hffffffff
)
)
===
1'bx
)
SVROKoIB
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRbONlu
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVROKoIB
!=
32'hffffffff
)
)
SVROKoIB
<=
SVROKoIB
+
32'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRGlDJE
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRGlDJE
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRGlDJE
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRUvXCJ
)
)
===
1'bx
)
SVRGlDJE
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRUvXCJ
)
)
SVRGlDJE
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRmNpYA
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRGlDJE
!=
32'hffffffff
)
)
===
1'bx
)
SVRGlDJE
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRmNpYA
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRGlDJE
!=
32'hffffffff
)
)
SVRGlDJE
<=
SVRGlDJE
+
32'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRczkkG
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRczkkG
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRczkkG
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRXKyOr
)
)
SVRczkkG
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRXKyOr
)
)
SVRczkkG
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRSMDrE
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRczkkG
!=
32'hffffffff
)
)
===
1'bx
)
SVRczkkG
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRSMDrE
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRczkkG
!=
32'hffffffff
)
)
SVRczkkG
<=
SVRczkkG
+
32'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRBmffQ
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRBmffQ
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRBmffQ
<=
32'd0
;
`ifdef SVRxoxPL 
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRKlIMZ
)
)
SVRBmffQ
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRKlIMZ
)
)
SVRBmffQ
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRwTOiP
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRBmffQ
!=
32'hffffffff
)
)
===
1'bx
)
SVRBmffQ
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRwTOiP
==
1'b1
)
&&
(
SVRnGCcv
==
1'b1
)
&&
(
SVRBmffQ
!=
32'hffffffff
)
)
SVRBmffQ
<=
SVRBmffQ
+
32'd1
;
assign
SVRoNaGz
=
SVRVyyGw
;
assign
SVRTmwId
=
SVRfJLFv
;
assign
SVRwglRb
=
SVROKoIB
;
assign
SVRxwbOR
=
SVRGlDJE
;
assign
SVRlLaUV
=
SVRczkkG
;
assign
SVRFsaXX
=
SVRBmffQ
;
endmodule
module SVRZiZDv
(
SVRJROZz
,
fclk
,
SVRrYaZV
,
SVRizAZX
,
SVRQfjSP
,
SVRhwAOL
,
SVRdlnUs
,
SVRBFgxj
)
;
input
SVRJROZz
;
input
fclk
;
input
[
23
:
0
]
SVRrYaZV
;
input
SVRizAZX
;
input
SVRQfjSP
;
input
SVRhwAOL
;
output
reg
[
23
:
0
]
SVRdlnUs
;
output
reg
SVRBFgxj
;
reg
[
15
:
0
]
SVRXpQwl
,
SVRYhvLf
;
reg
[
15
:
0
]
SVRlxgLT
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRXpQwl
<=
16'd640
;
SVRYhvLf
<=
16'd0
;
end
else
if
(
SVRQfjSP
==
1'b1
)
begin
SVRYhvLf
<=
16'd0
;
SVRXpQwl
<=
SVRYhvLf
;
end
else
if
(
SVRizAZX
==
1'b1
)
SVRYhvLf
<=
SVRYhvLf
+
16'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRlxgLT
<=
16'd0
;
else
if
(
SVRhwAOL
==
1'b1
)
SVRlxgLT
<=
16'd0
;
else
if
(
SVRQfjSP
==
1'b1
)
SVRlxgLT
<=
SVRlxgLT
+
16'd1
;
wire
[
15
:
0
]
SVRReZKN
=
SVRYhvLf
-
{
1'b0
,
SVRXpQwl
[
15
:
1
]
}
;
wire
[
3
:
0
]
SVRvCzSt
=
(
SVRXpQwl
>
2047
)
?
4'd8
:
(
SVRXpQwl
>
1024
)
?
4'd4
:
(
SVRXpQwl
>
512
)
?
4'd2
:
4'd1
;
wire
[
4
:
0
]
SVRwHIOa
=
(
SVRvCzSt
==
4'd1
)
?
SVRReZKN
[
4
:
0
]
:
(
SVRvCzSt
==
4'd2
)
?
SVRReZKN
[
5
:
1
]
:
(
SVRvCzSt
==
4'd4
)
?
SVRReZKN
[
6
:
2
]
:
SVRReZKN
[
7
:
3
]
;
wire
[
2
:
0
]
SVRXjNmR
=
(
SVRvCzSt
==
4'd1
)
?
SVRlxgLT
[
2
:
0
]
:
(
SVRvCzSt
==
4'd2
)
?
SVRlxgLT
[
3
:
1
]
:
(
SVRvCzSt
==
4'd4
)
?
SVRlxgLT
[
4
:
2
]
:
SVRlxgLT
[
5
:
3
]
;
wire
SVRkyPym
=
(
SVRReZKN
[
15
]
==
1'b1
)
?
1'b0
:
(
SVRReZKN
[
14
:
0
]
>
SVRvCzSt
*
32
)
?
1'b0
:
1'b1
;
wire
SVRrFQex
=
(
SVRlxgLT
>
8
*
SVRvCzSt
)
?
1'b0
:
1'b1
;
wire
SVRIpvCL
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd17
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd19
)
)
;
wire
SVRdBGGj
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRBnqQe
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRNgivc
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd23
)
||
(
SVRwHIOa
==
5'd24
)
||
(
SVRwHIOa
==
5'd25
)
||
(
SVRwHIOa
==
5'd26
)
||
(
SVRwHIOa
==
5'd27
)
)
;
wire
SVRtdEkB
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRJbpFn
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRdudIX
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd4
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd9
)
||
(
SVRwHIOa
==
5'd10
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd17
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd19
)
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRBFgxj
<=
1'd0
;
else
SVRBFgxj
<=
SVRizAZX
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRdlnUs
<=
24'd0
;
else
if
(
SVRkyPym
==
1'b0
)
SVRdlnUs
<=
SVRrYaZV
;
else
if
(
SVRrFQex
==
1'b0
)
SVRdlnUs
<=
SVRrYaZV
;
else
if
(
(
SVRXjNmR
==
3'd0
)
&&
(
SVRIpvCL
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd1
)
&&
(
SVRdBGGj
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd2
)
&&
(
SVRBnqQe
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd3
)
&&
(
SVRNgivc
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd4
)
&&
(
SVRtdEkB
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd5
)
&&
(
SVRJbpFn
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd6
)
&&
(
SVRdudIX
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
SVRdlnUs
<=
24'hFFFFFF
;
endmodule
module SVRwuuAu
(
SVRJROZz
,
fclk
,
SVRrYaZV
,
SVRizAZX
,
SVRQfjSP
,
SVRhwAOL
,
SVRdlnUs
,
SVRBFgxj
)
;
input
SVRJROZz
;
input
fclk
;
input
[
23
:
0
]
SVRrYaZV
;
input
SVRizAZX
;
input
SVRQfjSP
;
input
SVRhwAOL
;
output
reg
[
23
:
0
]
SVRdlnUs
;
output
reg
SVRBFgxj
;
reg
[
15
:
0
]
SVRXpQwl
,
SVRYhvLf
;
reg
[
15
:
0
]
SVRlxgLT
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRXpQwl
<=
16'd640
;
SVRYhvLf
<=
16'd0
;
end
else
if
(
SVRQfjSP
==
1'b1
)
begin
SVRYhvLf
<=
16'd0
;
SVRXpQwl
<=
SVRYhvLf
;
end
else
if
(
SVRizAZX
==
1'b1
)
SVRYhvLf
<=
SVRYhvLf
+
16'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRlxgLT
<=
16'd0
;
else
if
(
SVRhwAOL
==
1'b1
)
SVRlxgLT
<=
16'd0
;
else
if
(
SVRQfjSP
==
1'b1
)
SVRlxgLT
<=
SVRlxgLT
+
16'd1
;
wire
[
15
:
0
]
SVRReZKN
=
SVRYhvLf
-
{
1'b0
,
SVRXpQwl
[
15
:
1
]
}
;
wire
[
5
:
0
]
SVRvCzSt
=
(
SVRXpQwl
>
2047
)
?
6'd32
:
(
SVRXpQwl
>
1024
)
?
6'd16
:
(
SVRXpQwl
>
512
)
?
6'd8
:
4'd4
;
wire
[
4
:
0
]
SVRwHIOa
=
(
SVRvCzSt
==
6'd4
)
?
SVRReZKN
[
6
:
0
]
:
(
SVRvCzSt
==
6'd8
)
?
SVRReZKN
[
7
:
1
]
:
(
SVRvCzSt
==
6'd16
)
?
SVRReZKN
[
8
:
2
]
:
SVRReZKN
[
9
:
3
]
;
wire
[
2
:
0
]
SVRXjNmR
=
(
SVRvCzSt
==
6'd4
)
?
SVRlxgLT
[
4
:
0
]
:
(
SVRvCzSt
==
6'd8
)
?
SVRlxgLT
[
5
:
1
]
:
(
SVRvCzSt
==
6'd16
)
?
SVRlxgLT
[
6
:
2
]
:
SVRlxgLT
[
7
:
3
]
;
wire
SVRkyPym
=
(
SVRReZKN
[
15
]
==
1'b1
)
?
1'b0
:
(
SVRReZKN
[
14
:
0
]
>
SVRvCzSt
*
32
)
?
1'b0
:
1'b1
;
wire
SVRrFQex
=
1'b1
;
wire
SVRIpvCL
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd17
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd19
)
)
;
wire
SVRdBGGj
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRBnqQe
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRNgivc
=
(
(
SVRwHIOa
==
5'd2
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd6
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd23
)
||
(
SVRwHIOa
==
5'd24
)
||
(
SVRwHIOa
==
5'd25
)
||
(
SVRwHIOa
==
5'd26
)
||
(
SVRwHIOa
==
5'd27
)
)
;
wire
SVRtdEkB
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRJbpFn
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd5
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd12
)
||
(
SVRwHIOa
==
5'd15
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd25
)
)
;
wire
SVRdudIX
=
(
(
SVRwHIOa
==
5'd3
)
||
(
SVRwHIOa
==
5'd4
)
||
(
SVRwHIOa
==
5'd8
)
||
(
SVRwHIOa
==
5'd9
)
||
(
SVRwHIOa
==
5'd10
)
||
(
SVRwHIOa
==
5'd13
)
||
(
SVRwHIOa
==
5'd14
)
||
(
SVRwHIOa
==
5'd17
)
||
(
SVRwHIOa
==
5'd18
)
||
(
SVRwHIOa
==
5'd19
)
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRBFgxj
<=
1'd0
;
else
SVRBFgxj
<=
SVRizAZX
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRdlnUs
<=
24'd0
;
else
if
(
SVRkyPym
==
1'b0
)
SVRdlnUs
<=
SVRrYaZV
;
else
if
(
SVRrFQex
==
1'b0
)
SVRdlnUs
<=
SVRrYaZV
;
else
if
(
(
SVRXjNmR
==
3'd0
)
&&
(
SVRIpvCL
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd1
)
&&
(
SVRdBGGj
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd2
)
&&
(
SVRBnqQe
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd3
)
&&
(
SVRNgivc
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd4
)
&&
(
SVRtdEkB
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd5
)
&&
(
SVRJbpFn
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
if
(
(
SVRXjNmR
==
3'd6
)
&&
(
SVRdudIX
==
1'b1
)
)
SVRdlnUs
<=
24'd0
;
else
SVRdlnUs
<=
24'hFFFFFF
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRkYKaD
(
fclk
,
pclk
,
SVRyEtuR
,
SVRWiNOI
,
SVRzUTNy
,
SVRrGCzn
,
SVRehSHF
,
SVREusOH
,
SVRBdFMH
,
SVRCmjnh
,
SVRSCAjD
,
SVRgVTxt
,
SVRUtdgF
,
SVRHXUZw
,
SVRxZBBs
,
SVRXSjgA
,
SVRjDxvg
,
SVREOLkD
,
SVRBNOxF
,
SVRZmqEG
,
SVRoQJOJ
,
SVRAzazu
,
SVRklMnp
,
SVRbwSIu
,
SVRZfWeB
,
SVRTVbtZ
,
SVRZyNzG
,
SVRgDTYn
,
svr_fs
,
svr_fe
,
svr_ls
,
svr_le
,
svr_data_type
,
SVRoNaGz
,
SVRTmwId
,
SVRwglRb
,
SVRxwbOR
,
SVRlLaUV
,
SVRFsaXX
)
;
input
fclk
;
input
pclk
;
input
SVRyEtuR
;
input
SVRWiNOI
;
input
SVRzUTNy
;
input
SVRrGCzn
;
input
SVRehSHF
;
input
[
7
:
2
]
SVREusOH
;
input
[
7
:
2
]
SVRBdFMH
;
input
SVRCmjnh
;
input
SVRSCAjD
;
input
SVRgVTxt
;
input
wire
[
27
:
0
]
SVRUtdgF
;
input
wire
[
27
:
0
]
SVRHXUZw
;
`ifdef SVRsQYvh 
input
wire
[
31
:
0
]
SVRioKpl
;
`endif
input
wire
[
7
:
0
]
SVRxZBBs
;
input
wire
[
31
:
0
]
SVRXSjgA
;
input
wire
[
31
:
0
]
SVRjDxvg
;
input
wire
[
1
:
0
]
SVREOLkD
;
input
wire
[
31
:
0
]
SVRBNOxF
;
input
wire
[
31
:
0
]
SVRZmqEG
;
input
wire
SVRoQJOJ
;
input
wire
SVRAzazu
;
input
wire
[
7
:
0
]
SVRklMnp
;
input
wire
SVRbwSIu
;
input
wire
SVRZfWeB
;
output
[
31
:
0
]
SVRTVbtZ
;
output
wire
SVRZyNzG
;
output
reg
[
1
:
0
]
SVRgDTYn
;
output
reg
svr_fs
;
output
svr_fe
;
output
svr_ls
;
output
svr_le
;
`ifdef SVRyllEh 
output
SVRMFfPD
;
output
SVRTPCUO
;
`endif
output
reg
[
5
:
0
]
svr_data_type
;
`ifdef SVRNJLgb 
input
[
31
:
0
]
SVRoNaGz
;
input
[
31
:
0
]
SVRTmwId
;
input
[
31
:
0
]
SVRwglRb
;
input
[
31
:
0
]
SVRxwbOR
;
input
[
31
:
0
]
SVRlLaUV
;
input
[
31
:
0
]
SVRFsaXX
;
`endif
`ifdef SVRVOzuU 
input
[
31
:
0
]
SVRxUmkX
;
`endif
reg
SVRlxgFy
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRlxgFy
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVREusOH
,
2'b00
}
==
`SVRJyIko
)
)
===
1'bx
)
SVRlxgFy
<=
1'bx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVREusOH
,
2'b00
}
==
`SVRJyIko
)
)
SVRlxgFy
<=
SVRCmjnh
;
assign
SVRZyNzG
=
SVRlxgFy
;
wire
[
31
:
0
]
SVRReZhd
=
(
{
SVRBdFMH
,
2'b00
}
==
`SVRJyIko
)
?
{
31'd0
,
SVRlxgFy
}
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRDfNXx
)
?
{
4'd0
,
SVRUtdgF
}
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRawpRC
)
?
{
4'd0
,
SVRHXUZw
}
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRmEdoF
)
?
{
24'd0
,
SVRxZBBs
}
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRgPbHP
)
?
SVRXSjgA
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRPNWIl
)
?
SVRXSjgA
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRSfrTz
)
?
SVRjDxvg
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRWCIWM
)
?
SVREOLkD
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRyoryt
)
?
SVRBNOxF
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRmHiMj
)
?
SVRZmqEG
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRgnUJW
)
?
(
SVRgVTxt
)
?
SVRoNaGz
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRPZskp
)
?
(
SVRgVTxt
)
?
SVRTmwId
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRgtFxy
)
?
(
SVRgVTxt
)
?
SVRwglRb
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRUvXCJ
)
?
(
SVRgVTxt
)
?
SVRxwbOR
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRXKyOr
)
?
(
SVRgVTxt
)
?
SVRlLaUV
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRKlIMZ
)
?
(
SVRgVTxt
)
?
SVRFsaXX
:
32'd0
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRhnrhd
)
?
`SVRJNvGI
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRUqxEm
)
?
32'h00000206
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRJBHhX
)
?
32'h56_4C_53_49
:
(
{
SVRBdFMH
,
2'b00
}
==
`SVRRNQDy
)
?
32'h50_4C_55_53
:
32'h00000000
;
reg
[
31
:
0
]
SVRTVbtZ
;
always
@
(
posedge
pclk
or
negedge
SVRWiNOI
)
if
(
SVRWiNOI
==
1'b0
)
SVRTVbtZ
<=
32'h00000000
;
else
if
(
SVRrGCzn
&
~SVRSCAjD
&
SVRrGCzn
)
SVRTVbtZ
<=
SVRReZhd
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
svr_fs
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
svr_fs
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
svr_fs
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRklMnp
[
5
:
0
]
==
6'd0
)
&&
(
SVRbwSIu
==
1'b1
)
)
===
1'bx
)
svr_fs
<=
1'bx
;
`endif
else
if
(
(
SVRklMnp
[
5
:
0
]
==
6'd0
)
&&
(
SVRbwSIu
==
1'b1
)
)
svr_fs
<=
1'b1
;
else
svr_fs
<=
1'b0
;
reg
SVRvCZDB
;
reg
SVRwHvHE
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRvCZDB
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRvCZDB
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRvCZDB
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRbwSIu
&
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
&
~SVRwHvHE
)
===
1'bx
)
SVRvCZDB
<=
1'bx
;
`endif
else
if
(
SVRbwSIu
&
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
&
~SVRwHvHE
)
SVRvCZDB
<=
1'b1
;
else
SVRvCZDB
<=
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRwHvHE
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRwHvHE
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRwHvHE
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRbwSIu
&
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
)
===
1'bx
)
SVRwHvHE
<=
1'bx
;
`endif
else
if
(
SVRbwSIu
&
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
)
SVRwHvHE
<=
1'b1
;
else
SVRwHvHE
<=
1'b0
;
assign
svr_fe
=
SVRvCZDB
;
reg
[
1
:
0
]
SVRXJgjG
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRXJgjG
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
SVRZfWeB
===
1'bx
)
SVRXJgjG
<=
2'bxx
;
`endif
else
if
(
SVRZfWeB
)
SVRXJgjG
<=
2'b01
;
else
SVRXJgjG
<=
{
SVRXJgjG
[
0
]
,
1'b0
}
;
assign
svr_ls
=
(
SVRXJgjG
!=
2'b01
)
?
1'b0
:
1'b1
;
reg
SVRYrDeq
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRYrDeq
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRoQJOJ
)
===
1'bx
)
SVRYrDeq
<=
1'bx
;
`endif
else
if
(
(
SVRoQJOJ
)
)
SVRYrDeq
<=
1'b1
;
else
SVRYrDeq
<=
1'b0
;
assign
svr_le
=
(
SVRYrDeq
)
?
1'b0
:
(
SVRoQJOJ
)
?
1'b1
:
1'b0
;
`ifdef SVRyllEh 
reg
SVRZIoci
,
SVRzrhbE
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRZIoci
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd2
)
)
===
1'bx
)
SVRZIoci
<=
1'bx
;
`endif
else
if
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd2
)
)
SVRZIoci
<=
1'b1
;
else
SVRZIoci
<=
1'b0
;
assign
SVRMFfPD
=
(
SVRZIoci
==
1'b1
)
?
1'b0
:
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd2
)
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRzrhbE
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd3
)
)
===
1'bx
)
SVRzrhbE
<=
1'bx
;
`endif
else
if
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd3
)
)
SVRzrhbE
<=
1'b1
;
else
SVRzrhbE
<=
1'b0
;
assign
SVRTPCUO
=
(
SVRzrhbE
==
1'b1
)
?
1'b0
:
(
(
SVRbwSIu
)
&&
(
SVRklMnp
[
5
:
0
]
==
6'd3
)
)
?
1'b1
:
1'b0
;
`endif
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRgDTYn
<=
2'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRgDTYn
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRgDTYn
<=
2'd0
;
else
SVRgDTYn
<=
SVRklMnp
[
7
:
6
]
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
svr_data_type
<=
6'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
svr_data_type
<=
6'bxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
svr_data_type
<=
6'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRbwSIu
==
1'b1
)
===
1'bx
)
svr_data_type
<=
6'bxx_xxxx
;
`endif
else
if
(
SVRbwSIu
==
1'b1
)
svr_data_type
<=
SVRklMnp
[
5
:
0
]
;
endmodule
module SVRBMFcH
(
SVRaPJKf
,
SVRyMoCu
,
SVRDXWLJ
,
SVRasuLi
,
SVRmcglv
,
SVRmthok
,
SVRSCzZV
,
SVRIHiSO
)
;
input
SVRaPJKf
;
input
[
31
:
0
]
SVRyMoCu
;
input
[
31
:
0
]
SVRDXWLJ
;
input
[
31
:
0
]
SVRasuLi
;
input
[
31
:
0
]
SVRmcglv
;
output
SVRmthok
;
output
SVRSCzZV
;
output
SVRIHiSO
;
localparam
SVRMIDap
=
32'h5648FEB3
;
localparam
SVRFKKsY
=
32'hEE687CE6
;
localparam
SVRpssjz
=
32'h046E11EA
;
localparam
SVRtcfxD
=
32'hC09A1BB4
;
localparam
SVRjBCLO
=
32'h0C7D1DDA
;
localparam
SVRQgklL
=
32'hF7F3E9FC
;
localparam
SVRvdFFS
=
32'h1E250431
;
localparam
SVRWuliN
=
32'h21B55210
;
localparam
SVRyKfET
=
32'hF879CFEB
;
localparam
SVRyLyHN
=
32'h662E1359
;
localparam
SVRYliJK
=
32'h76318F1E
;
localparam
SVRlZZjj
=
32'hD9DA5DD1
;
localparam
SVRRSvxv
=
32'h67C14A63
;
localparam
SVRvWKLK
=
32'hA2BF06C2
;
localparam
SVRwrolj
=
32'h7DE71358
;
wire
[
31
:
0
]
SVRXbdyV
,
SVRkuxEo
,
SVRrDHhy
,
SVRUHmWC
,
SVRXqgyO
;
wire
[
31
:
0
]
SVRKbzel
,
SVReuIuW
,
SVRckrky
,
SVRnyEXc
,
SVRgmPyb
;
wire
[
31
:
0
]
SVRdGuMa
,
SVRnjGlr
,
SVRSXlyz
,
SVRWYfMm
,
SVRKSylX
;
assign
SVRXbdyV
=
SVRyMoCu
^
SVRMIDap
;
assign
SVRKbzel
=
SVRyMoCu
^
SVRFKKsY
;
assign
SVRdGuMa
=
SVRyMoCu
^
SVRpssjz
;
SVRswMFY
SVRvepiQ
(
SVRaPJKf
,
SVRXbdyV
,
SVRtcfxD
,
SVRkuxEo
)
;
SVRswMFY
SVRwvDWL
(
SVRaPJKf
,
SVRKbzel
,
SVRjBCLO
,
SVReuIuW
)
;
SVRswMFY
SVRXDKQj
(
SVRaPJKf
,
SVRdGuMa
,
SVRQgklL
,
SVRnjGlr
)
;
SVRswMFY
SVRkiONv
(
SVRaPJKf
,
SVRkuxEo
,
SVRvdFFS
,
SVRrDHhy
)
;
SVRswMFY
SVRrXpMB
(
SVRaPJKf
,
SVReuIuW
,
SVRWuliN
,
SVRckrky
)
;
SVRswMFY
SVRURDLE
(
SVRaPJKf
,
SVRnjGlr
,
SVRyKfET
,
SVRSXlyz
)
;
SVRswMFY
SVRjPklG
(
SVRaPJKf
,
SVRrDHhy
,
SVRyLyHN
,
SVRUHmWC
)
;
SVRswMFY
SVREuFfQ
(
SVRaPJKf
,
SVRckrky
,
SVRYliJK
,
SVRnyEXc
)
;
SVRswMFY
SVRBDlVl
(
SVRaPJKf
,
SVRSXlyz
,
SVRlZZjj
,
SVRWYfMm
)
;
SVRswMFY
SVRNOFXf
(
SVRaPJKf
,
SVRUHmWC
,
SVRRSvxv
,
SVRXqgyO
)
;
SVRswMFY
SVRFNlRT
(
SVRaPJKf
,
SVRnyEXc
,
SVRvWKLK
,
SVRgmPyb
)
;
SVRswMFY
SVRPTFVW
(
SVRaPJKf
,
SVRWYfMm
,
SVRwrolj
,
SVRKSylX
)
;
reg
SVRmthok
,
SVRSCzZV
,
SVRIHiSO
;
initial
SVRmthok
=
1'b0
;
initial
SVRSCzZV
=
1'b0
;
initial
SVRIHiSO
=
1'b0
;
always
@
(
posedge
SVRaPJKf
)
if
(
SVRXqgyO
==
SVRDXWLJ
)
SVRmthok
<=
1'b1
;
else
SVRmthok
<=
1'b0
;
always
@
(
posedge
SVRaPJKf
)
if
(
SVRgmPyb
==
SVRasuLi
)
SVRSCzZV
<=
1'b1
;
else
SVRSCzZV
<=
1'b0
;
always
@
(
posedge
SVRaPJKf
)
if
(
SVRKSylX
==
SVRmcglv
)
SVRIHiSO
<=
1'b1
;
else
SVRIHiSO
<=
1'b0
;
endmodule
module SVRswMFY
(
SVRaPJKf
,
SVRAopDX
,
SVRvovDu
,
SVRUWPxY
)
;
input
SVRaPJKf
;
input
[
31
:
0
]
SVRAopDX
;
input
[
31
:
0
]
SVRvovDu
;
output
[
31
:
0
]
SVRUWPxY
;
wire
[
31
:
0
]
SVRJRqeq
,
SVRRvicI
,
SVRVkebR
,
SVRJYXsm
,
SVRrZyjG
,
SVRIzMeQ
;
SVRRmtcv
SVRvGjBk
(
SVRAopDX
,
SVRvovDu
[
4
:
0
]
,
SVRJRqeq
)
;
SVRRmtcv
SVRwJagW
(
SVRJRqeq
,
SVRvovDu
[
9
:
5
]
,
SVRRvicI
)
;
SVRRmtcv
SVRLrady
(
SVRRvicI
,
SVRvovDu
[
14
:
10
]
,
SVRVkebR
)
;
SVRRmtcv
SVRSiAbM
(
SVRVkebR
,
SVRvovDu
[
19
:
15
]
,
SVRJYXsm
)
;
SVRRmtcv
SVRIXiTj
(
SVRJYXsm
,
SVRvovDu
[
24
:
20
]
,
SVRrZyjG
)
;
SVRRmtcv
SVRRyEWE
(
SVRrZyjG
,
SVRvovDu
[
29
:
25
]
,
SVRIzMeQ
)
;
reg
[
7
:
0
]
SVRvmpyP
,
SVRwzDEl
,
SVRXFKHw
,
SVRYpSql
;
always
@
(
posedge
SVRaPJKf
)
case
(
SVRvovDu
[
31
:
30
]
)
2'b00
:
begin
SVRvmpyP
<=
SVRIzMeQ
[
15
:
8
]
;
SVRwzDEl
<=
SVRIzMeQ
[
7
:
0
]
;
SVRXFKHw
<=
SVRIzMeQ
[
31
:
24
]
;
SVRYpSql
<=
SVRIzMeQ
[
23
:
16
]
;
end
2'b01
:
begin
SVRvmpyP
<=
SVRIzMeQ
[
23
:
16
]
;
SVRwzDEl
<=
SVRIzMeQ
[
31
:
24
]
;
SVRXFKHw
<=
SVRIzMeQ
[
7
:
0
]
;
SVRYpSql
<=
SVRIzMeQ
[
15
:
8
]
;
end
2'b10
:
begin
SVRvmpyP
<=
SVRIzMeQ
[
15
:
8
]
;
SVRwzDEl
<=
SVRIzMeQ
[
23
:
16
]
;
SVRXFKHw
<=
SVRIzMeQ
[
31
:
24
]
;
SVRYpSql
<=
SVRIzMeQ
[
7
:
0
]
;
end
2'b11
:
begin
SVRvmpyP
<=
SVRIzMeQ
[
31
:
24
]
;
SVRwzDEl
<=
SVRIzMeQ
[
7
:
0
]
;
SVRXFKHw
<=
SVRIzMeQ
[
15
:
8
]
;
SVRYpSql
<=
SVRIzMeQ
[
23
:
16
]
;
end
default
:
begin
SVRvmpyP
<=
8'd0
;
SVRwzDEl
<=
8'd0
;
SVRXFKHw
<=
8'd0
;
SVRYpSql
<=
8'd0
;
end
endcase
assign
SVRUWPxY
=
{
SVRYpSql
,
SVRXFKHw
,
SVRwzDEl
,
SVRvmpyP
}
;
endmodule
module SVRRmtcv
(
SVRAopDX
,
SVRvovDu
,
SVRUWPxY
)
;
input
[
31
:
0
]
SVRAopDX
;
input
[
4
:
0
]
SVRvovDu
;
output
[
31
:
0
]
SVRUWPxY
;
wire
SVRlbSAW
=
SVRAopDX
[
SVRvovDu
]
;
wire
[
31
:
0
]
SVRFawnY
=
(
SVRvovDu
==
5'd
0
)
?
32'h00000001
:
(
SVRvovDu
==
5'd
1
)
?
32'h00000002
:
(
SVRvovDu
==
5'd
2
)
?
32'h00000004
:
(
SVRvovDu
==
5'd
3
)
?
32'h00000008
:
(
SVRvovDu
==
5'd
4
)
?
32'h00000010
:
(
SVRvovDu
==
5'd
5
)
?
32'h00000020
:
(
SVRvovDu
==
5'd
6
)
?
32'h00000040
:
(
SVRvovDu
==
5'd
7
)
?
32'h00000080
:
(
SVRvovDu
==
5'd
8
)
?
32'h00000100
:
(
SVRvovDu
==
5'd
9
)
?
32'h00000200
:
(
SVRvovDu
==
5'd10
)
?
32'h00000400
:
(
SVRvovDu
==
5'd11
)
?
32'h00000800
:
(
SVRvovDu
==
5'd12
)
?
32'h00001000
:
(
SVRvovDu
==
5'd13
)
?
32'h00002000
:
(
SVRvovDu
==
5'd14
)
?
32'h00004000
:
(
SVRvovDu
==
5'd15
)
?
32'h00008000
:
(
SVRvovDu
==
5'd16
)
?
32'h00010000
:
(
SVRvovDu
==
5'd17
)
?
32'h00020000
:
(
SVRvovDu
==
5'd18
)
?
32'h00040000
:
(
SVRvovDu
==
5'd19
)
?
32'h00080000
:
(
SVRvovDu
==
5'd20
)
?
32'h00100000
:
(
SVRvovDu
==
5'd21
)
?
32'h00200000
:
(
SVRvovDu
==
5'd22
)
?
32'h00400000
:
(
SVRvovDu
==
5'd23
)
?
32'h00800000
:
(
SVRvovDu
==
5'd24
)
?
32'h01000000
:
(
SVRvovDu
==
5'd25
)
?
32'h02000000
:
(
SVRvovDu
==
5'd26
)
?
32'h04000000
:
(
SVRvovDu
==
5'd27
)
?
32'h08000000
:
(
SVRvovDu
==
5'd28
)
?
32'h10000000
:
(
SVRvovDu
==
5'd29
)
?
32'h20000000
:
(
SVRvovDu
==
5'd30
)
?
32'h40000000
:
32'h80000000
;
assign
SVRUWPxY
=
(
SVRvovDu
==
5'd0
)
?
SVRAopDX
:
(
SVRAopDX
[
0
]
==
1'b0
)
?
{
SVRAopDX
[
31
:
1
]
,
SVRlbSAW
}
&
~SVRFawnY
:
{
SVRAopDX
[
31
:
1
]
,
SVRlbSAW
}
|
SVRFawnY
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRZuLLH
(
fclk
,
SVRJROZz
,
SVRehSHF
,
SVRyMsqX
,
SVRmtjIy
,
SVRUtdgF
,
SVRHXUZw
,
SVRSoHSD
,
SVRwHqWo
,
SVRXjEqy
)
;
input
wire
fclk
;
input
wire
SVRJROZz
;
input
wire
SVRehSHF
;
input
wire
[
7
:
2
]
SVRyMsqX
;
input
wire
[
31
:
0
]
SVRmtjIy
;
output
[
27
:
0
]
SVRUtdgF
;
output
[
27
:
0
]
SVRHXUZw
;
output
[
31
:
0
]
SVRSoHSD
;
output
[
31
:
0
]
SVRwHqWo
;
output
[
31
:
0
]
SVRXjEqy
;
reg
[
27
:
0
]
SVRntUoD
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRntUoD
<=
28'd11 // 9-April-2015 change (was 28'd1)
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRDfNXx
)
)
===
1'bx
)
SVRntUoD
<=
28'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRDfNXx
)
)
SVRntUoD
<=
SVRmtjIy
[
27
:
0
]
;
reg
[
27
:
0
]
SVRGjxHo
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRGjxHo
<=
28'h0000000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRawpRC
)
)
===
1'bx
)
SVRGjxHo
<=
28'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRawpRC
)
)
SVRGjxHo
<=
{
~SVRmtjIy
[
27
:
24
]
,
SVRmtjIy
[
23
:
0
]
}
;
reg
[
31
:
0
]
SVRQELqH
;
always
@
(
posedge
fclk
)
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRDGIDb
)
)
SVRQELqH
<=
SVRmtjIy
;
reg
[
31
:
0
]
SVRvPsIq
;
always
@
(
posedge
fclk
)
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRoqROa
)
)
SVRvPsIq
<=
SVRmtjIy
;
reg
[
31
:
0
]
SVRKujri
;
always
@
(
posedge
fclk
)
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRtBRmr
)
)
SVRKujri
<=
SVRmtjIy
;
initial
#
0
begin
SVRQELqH
=
32'd0
;
SVRvPsIq
=
32'd0
;
SVRKujri
=
32'd0
;
end
assign
SVRSoHSD
=
SVRQELqH
;
assign
SVRwHqWo
=
SVRvPsIq
;
assign
SVRXjEqy
=
SVRKujri
;
assign
SVRUtdgF
=
SVRntUoD
;
assign
SVRHXUZw
=
{
~SVRGjxHo
[
27
:
24
]
,
SVRGjxHo
[
23
:
0
]
}
;
`ifdef	PROG_CSI_SYNC
reg
[
31
:
0
]
SVRsKEie
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRsKEie
<=
32'hb8b8b8b8
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRqiCwc
)
)
===
1'bx
)
SVRsKEie
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRqiCwc
)
)
SVRsKEie
<=
SVRmtjIy
;
assign
SVRioKpl
=
SVRsKEie
;
`endif
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
`define SVRPyLMf            6'h10
`define SVRuMsTc         3'b010
`define SVRwmfpS          6'h1A
`define SVRlGChw          6'b011000
`define SVRfqOdL          6'b011100
`define SVRobquj         6'b011001
`define SVRHaiKE         6'b011101
`define SVRCTzkG           6'b01_1110
`define SVROWmfQ          6'b01_1111
`define SVRGrcVL          6'b10_0000
`define SVRQiBXS          6'b10_0001
`define SVRHxjrN          6'b10_0010
`define SVRQLEIT          6'b10_0011
`define SVRhmLJN          6'b10_0100
`define SVRpzoKK            6'b10_1000
`define SVRTfDkj            6'b10_1001
`define SVRiwKxv            6'b10_1010
`define SVRelSLK           6'b10_1011
`define SVRCfWss           6'b10_1100
`define SVROcyjJ           6'b10_1101
`define SVRubMEr             6'b11_0000
module SVRFoNQp
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRknrFe
,
SVRsUANj
,
SVRoAAnA
,
SVRVmcEw
,
SVRGKeQn
,
SVRxgbpl
,
SVRoQJOJ
,
SVRBcWQp
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRzUTNy
;
input
[
15
:
0
]
SVRknrFe
;
input
SVRsUANj
;
input
SVRoAAnA
;
output
[
23
:
0
]
SVRVmcEw
;
input
[
5
:
0
]
SVRGKeQn
;
output
SVRxgbpl
;
output
SVRoQJOJ
;
input
SVRBcWQp
;
wire
SVRWTOHZ
;
wire
[
3
:
0
]
SVRYwUQz
,
SVRLeTND
;
wire
[
9
:
0
]
SVREvsMF
;
wire
[
3
:
0
]
SVRPkjTp
=
(
SVRGKeQn
==
`SVRPyLMf
)
?
4'h0
:
(
SVRGKeQn
[
5
:
3
]
==
`SVRuMsTc
)
?
4'h0
:
(
SVRGKeQn
==
`SVRwmfpS
)
?
4'h0
:
(
SVRGKeQn
==
`SVRlGChw
)
?
4'h0
:
(
SVRGKeQn
==
`SVRfqOdL
)
?
4'h0
:
(
SVRGKeQn
==
`SVRCTzkG
)
?
4'h0
:
(
SVRGKeQn
==
`SVRiwKxv
)
?
4'h0
:
(
SVRGKeQn
==
`SVRubMEr
)
?
4'h0
:
(
SVRGKeQn
==
`SVRelSLK
)
?
4'h1
:
(
SVRGKeQn
==
`SVRCfWss
)
?
4'ha
:
(
SVRGKeQn
==
`SVROWmfQ
)
?
4'h1
:
(
SVRGKeQn
==
`SVRobquj
)
?
4'h1
:
(
SVRGKeQn
==
`SVRHaiKE
)
?
4'h1
:
(
SVRGKeQn
==
`SVRGrcVL
)
?
4'h2
:
(
SVRGKeQn
==
`SVRQiBXS
)
?
4'h3
:
(
SVRGKeQn
==
`SVRHxjrN
)
?
4'h4
:
(
SVRGKeQn
==
`SVRQLEIT
)
?
4'h5
:
(
SVRGKeQn
==
`SVRhmLJN
)
?
4'h6
:
(
SVRGKeQn
==
`SVRpzoKK
)
?
4'h7
:
(
SVRGKeQn
==
`SVRTfDkj
)
?
4'h8
:
(
SVRGKeQn
==
`SVRelSLK
)
?
4'h1
:
(
SVRGKeQn
==
`SVRCfWss
)
?
4'ha
:
(
SVRGKeQn
==
`SVROcyjJ
)
?
4'hb
:
4'h0
;
reg
[
15
:
0
]
SVRGyaPY
[
4
:
0
]
;
reg
[
2
:
0
]
SVRqmAuZ
;
reg
[
3
:
0
]
SVRignKZ
;
reg
SVReDgSz
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVReDgSz
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVReDgSz
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVReDgSz
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVReDgSz
==
1'b0
)
&&
(
SVRoAAnA
==
1'b1
)
)
===
1'bx
)
SVReDgSz
<=
1'bx
;
`endif
else
if
(
(
SVReDgSz
==
1'b0
)
&&
(
SVRoAAnA
==
1'b1
)
)
SVReDgSz
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVREvsMF
[
2
]
==
1'b0
)
&&
(
SVRoAAnA
==
1'b0
)
)
===
1'bx
)
SVReDgSz
<=
1'bx
;
`endif
else
if
(
(
SVREvsMF
[
2
]
==
1'b0
)
&&
(
SVRoAAnA
==
1'b0
)
)
SVReDgSz
<=
1'b0
;
wire
SVROhzOd
=
SVRoAAnA
|
SVReDgSz
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRGyaPY
[
0
]
<=
16'd0
;
SVRGyaPY
[
1
]
<=
16'd0
;
SVRGyaPY
[
2
]
<=
16'd0
;
SVRGyaPY
[
3
]
<=
16'd0
;
SVRGyaPY
[
4
]
<=
16'd0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRsUANj
==
1'b1
)
===
1'bx
)
SVRGyaPY
[
SVRqmAuZ
]
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRsUANj
==
1'b1
)
SVRGyaPY
[
SVRqmAuZ
]
<=
SVRknrFe
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRqmAuZ
<=
3'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVROhzOd
==
1'b0
)
===
1'bx
)
SVRqmAuZ
<=
3'bxxx
;
`endif
else
if
(
SVROhzOd
==
1'b0
)
SVRqmAuZ
<=
3'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRsUANj
==
1'b1
)
&&
(
SVRqmAuZ
==
3'd4
)
)
===
1'bx
)
SVRqmAuZ
<=
3'bxxx
;
`endif
else
if
(
(
SVRsUANj
==
1'b1
)
&&
(
SVRqmAuZ
==
3'd4
)
)
SVRqmAuZ
<=
3'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRsUANj
==
1'b1
)
===
1'bx
)
SVRqmAuZ
<=
3'bxxx
;
`endif
else
if
(
SVRsUANj
==
1'b1
)
SVRqmAuZ
<=
SVRqmAuZ
+
3'd1
;
wire
[
9
:
0
]
SVRUDmUB
=
(
(
SVRBcWQp
==
1'b0
)
&&
(
SVRqmAuZ
==
3'b000
)
)
?
10'b0000000011
:
(
(
SVRBcWQp
==
1'b0
)
&&
(
SVRqmAuZ
==
3'b001
)
)
?
10'b0000001100
:
(
(
SVRBcWQp
==
1'b0
)
&&
(
SVRqmAuZ
==
3'b010
)
)
?
10'b0000110000
:
(
(
SVRBcWQp
==
1'b0
)
&&
(
SVRqmAuZ
==
3'b011
)
)
?
10'b0011000000
:
(
(
SVRBcWQp
==
1'b0
)
&&
(
SVRqmAuZ
==
3'b100
)
)
?
10'b1100000000
:
(
(
SVRBcWQp
==
1'b1
)
&&
(
SVRqmAuZ
==
3'b000
)
)
?
10'b0000000001
:
(
(
SVRBcWQp
==
1'b1
)
&&
(
SVRqmAuZ
==
3'b001
)
)
?
10'b0000000100
:
(
(
SVRBcWQp
==
1'b1
)
&&
(
SVRqmAuZ
==
3'b010
)
)
?
10'b0000010000
:
(
(
SVRBcWQp
==
1'b1
)
&&
(
SVRqmAuZ
==
3'b011
)
)
?
10'b0001000000
:
10'b0100000000
;
wire
[
3
:
0
]
SVRXogXN
=
(
SVRPkjTp
==
4'h0
)
?
4'd1
:
(
SVRPkjTp
==
4'h1
)
?
4'd5
:
(
SVRPkjTp
==
4'h2
)
?
4'd2
:
(
SVRPkjTp
==
4'h3
)
?
4'd2
:
(
SVRPkjTp
==
4'h4
)
?
4'd2
:
(
SVRPkjTp
==
4'h5
)
?
4'd9
:
(
SVRPkjTp
==
4'h6
)
?
4'd3
:
(
SVRPkjTp
==
4'h7
)
?
4'd3
:
(
SVRPkjTp
==
4'h8
)
?
4'd7
:
(
SVRPkjTp
==
4'ha
)
?
4'd3
:
(
SVRPkjTp
==
4'hb
)
?
4'd7
:
4'd1
;
wire
[
9
:
0
]
SVRyhDYt
=
(
SVRXogXN
==
4'b0001
)
?
10'b0000000001
:
(
SVRXogXN
==
4'b0010
)
?
10'b0000000011
:
(
SVRXogXN
==
4'b0011
)
?
10'b0000000111
:
(
SVRXogXN
==
4'b0100
)
?
10'b0000001111
:
(
SVRXogXN
==
4'b0101
)
?
10'b0000011111
:
(
SVRXogXN
==
4'b0110
)
?
10'b0000111111
:
(
SVRXogXN
==
4'b0111
)
?
10'b0001111111
:
(
SVRXogXN
==
4'b1000
)
?
10'b0011111111
:
10'b0111111111
;
wire
[
9
:
0
]
SVRMDoZj
=
(
SVRignKZ
==
4'b0000
)
?
{
SVRyhDYt
}
:
(
SVRignKZ
==
4'b0001
)
?
{
SVRyhDYt
[
8
:
0
]
,
SVRyhDYt
[
9
]
}
:
(
SVRignKZ
==
4'b0010
)
?
{
SVRyhDYt
[
7
:
0
]
,
SVRyhDYt
[
9
:
8
]
}
:
(
SVRignKZ
==
4'b0011
)
?
{
SVRyhDYt
[
6
:
0
]
,
SVRyhDYt
[
9
:
7
]
}
:
(
SVRignKZ
==
4'b0100
)
?
{
SVRyhDYt
[
5
:
0
]
,
SVRyhDYt
[
9
:
6
]
}
:
(
SVRignKZ
==
4'b0101
)
?
{
SVRyhDYt
[
4
:
0
]
,
SVRyhDYt
[
9
:
5
]
}
:
(
SVRignKZ
==
4'b0110
)
?
{
SVRyhDYt
[
3
:
0
]
,
SVRyhDYt
[
9
:
4
]
}
:
(
SVRignKZ
==
4'b0111
)
?
{
SVRyhDYt
[
2
:
0
]
,
SVRyhDYt
[
9
:
3
]
}
:
(
SVRignKZ
==
4'b1000
)
?
{
SVRyhDYt
[
1
:
0
]
,
SVRyhDYt
[
9
:
2
]
}
:
{
SVRyhDYt
[
0
]
,
SVRyhDYt
[
9
:
1
]
}
;
reg
[
9
:
0
]
SVRfidSV
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRfidSV
<=
10'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVROhzOd
==
1'b0
)
===
1'bx
)
SVRfidSV
<=
10'bxx_xxxx_xxxx
;
`endif
else
if
(
SVROhzOd
==
1'b0
)
SVRfidSV
<=
10'd0
;
else
SVRfidSV
<=
(
SVRUDmUB
&
{
10
{
SVRoAAnA
}
}
&
{
10
{
SVRsUANj
}
}
)
|
(
SVRfidSV
&
~
(
SVRMDoZj
&
{
10
{
SVRWTOHZ
}
}
)
)
;
wire
[
4
:
0
]
SVRoxxOo
=
(
{
1'b0
,
SVRignKZ
}
+
{
1'b0
,
SVRLeTND
}
)
;
wire
[
4
:
0
]
SVRTEHmY
=
(
SVRoxxOo
-
5'd10
)
;
wire
[
3
:
0
]
SVRIIMYp
=
(
SVRoxxOo
>=
5'd10
)
?
SVRTEHmY
[
3
:
0
]
:
SVRoxxOo
[
3
:
0
]
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRignKZ
<=
4'd0
;
else
if
(
SVRzUTNy
==
1'b1
)
SVRignKZ
<=
4'd0
;
else
if
(
~SVROhzOd
)
SVRignKZ
<=
4'd0
;
else
if
(
SVRWTOHZ
)
SVRignKZ
<=
SVRIIMYp
;
wire
[
71
:
0
]
SVRDkPRy
=
(
SVRignKZ
==
4'b0000
)
?
{
SVRGyaPY
[
4
]
[
7
:
0
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
}
:
(
SVRignKZ
==
4'b0001
)
?
{
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
[
15
:
8
]
}
:
(
SVRignKZ
==
4'b0010
)
?
{
SVRGyaPY
[
0
]
[
7
:
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
}
:
(
SVRignKZ
==
4'b0011
)
?
{
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
[
15
:
8
]
}
:
(
SVRignKZ
==
4'b0100
)
?
{
SVRGyaPY
[
1
]
[
7
:
0
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
}
:
(
SVRignKZ
==
4'b0101
)
?
{
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
[
15
:
8
]
}
:
(
SVRignKZ
==
4'b0110
)
?
{
SVRGyaPY
[
2
]
[
7
:
0
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
}
:
(
SVRignKZ
==
4'b0111
)
?
{
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
,
SVRGyaPY
[
3
]
[
15
:
8
]
}
:
(
SVRignKZ
==
4'b1000
)
?
{
SVRGyaPY
[
3
]
[
7
:
0
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
}
:
{
SVRGyaPY
[
3
]
,
SVRGyaPY
[
2
]
,
SVRGyaPY
[
1
]
,
SVRGyaPY
[
0
]
,
SVRGyaPY
[
4
]
[
15
:
8
]
}
;
assign
SVREvsMF
=
(
SVRignKZ
==
4'b0000
)
?
SVRfidSV
:
(
SVRignKZ
==
4'b0001
)
?
{
SVRfidSV
[
0
]
,
SVRfidSV
[
9
:
1
]
}
:
(
SVRignKZ
==
4'b0010
)
?
{
SVRfidSV
[
1
:
0
]
,
SVRfidSV
[
9
:
2
]
}
:
(
SVRignKZ
==
4'b0011
)
?
{
SVRfidSV
[
2
:
0
]
,
SVRfidSV
[
9
:
3
]
}
:
(
SVRignKZ
==
4'b0100
)
?
{
SVRfidSV
[
3
:
0
]
,
SVRfidSV
[
9
:
4
]
}
:
(
SVRignKZ
==
4'b0101
)
?
{
SVRfidSV
[
4
:
0
]
,
SVRfidSV
[
9
:
5
]
}
:
(
SVRignKZ
==
4'b0110
)
?
{
SVRfidSV
[
5
:
0
]
,
SVRfidSV
[
9
:
6
]
}
:
(
SVRignKZ
==
4'b0111
)
?
{
SVRfidSV
[
6
:
0
]
,
SVRfidSV
[
9
:
7
]
}
:
(
SVRignKZ
==
4'b1000
)
?
{
SVRfidSV
[
7
:
0
]
,
SVRfidSV
[
9
:
8
]
}
:
{
SVRfidSV
[
8
:
0
]
,
SVRfidSV
[
9
]
}
;
wire
SVRAyqoD
=
(
(
SVRXogXN
==
4'b0001
)
&&
(
SVREvsMF
[
0
]
==
1'b1
)
)
?
1'b1
:
(
(
SVRXogXN
==
4'b0010
)
&&
(
SVREvsMF
[
1
]
==
1'b1
)
)
?
1'b1
:
(
(
SVRXogXN
==
4'b0011
)
&&
(
SVREvsMF
[
2
]
==
1'b1
)
)
?
1'b1
:
(
(
SVRXogXN
==
4'b0101
)
&&
(
SVREvsMF
[
4
]
==
1'b1
)
)
?
1'b1
:
(
(
SVRXogXN
==
4'b0111
)
&&
(
SVREvsMF
[
6
]
==
1'b1
)
)
?
1'b1
:
(
(
SVRXogXN
==
4'b1001
)
&&
(
SVREvsMF
[
8
]
==
1'b1
)
)
?
1'b1
:
1'b0
;
wire
SVRzfEzF
;
assign
SVRWTOHZ
=
(
SVRAyqoD
&
SVRzfEzF
)
;
reg
[
71
:
0
]
SVRMcPMP
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRMcPMP
<=
72'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRWTOHZ
)
===
1'bx
)
SVRMcPMP
<=
80'bxxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx_xxxxxxxx
;
`endif
else
if
(
SVRWTOHZ
)
SVRMcPMP
<=
SVRDkPRy
;
assign
SVRYwUQz
=
(
SVRPkjTp
==
4'h0
)
?
4'd1
:
(
SVRPkjTp
==
4'h1
)
?
4'd4
:
(
SVRPkjTp
==
4'h2
)
?
4'd1
:
(
SVRPkjTp
==
4'h3
)
?
4'd1
:
(
SVRPkjTp
==
4'h4
)
?
4'd1
:
(
SVRPkjTp
==
4'h5
)
?
4'd4
:
(
SVRPkjTp
==
4'h6
)
?
4'd1
:
(
SVRPkjTp
==
4'h7
)
?
4'd4
:
(
SVRPkjTp
==
4'h8
)
?
4'd8
:
(
SVRPkjTp
==
4'ha
)
?
4'd2
:
(
SVRPkjTp
==
4'hb
)
?
4'd4
:
4'd0
;
assign
SVRLeTND
=
(
SVRPkjTp
==
4'h0
)
?
4'd1
:
(
SVRPkjTp
==
4'h1
)
?
4'd5
:
(
SVRPkjTp
==
4'h2
)
?
4'd2
:
(
SVRPkjTp
==
4'h3
)
?
4'd2
:
(
SVRPkjTp
==
4'h4
)
?
4'd2
:
(
SVRPkjTp
==
4'h5
)
?
4'd9
:
(
SVRPkjTp
==
4'h6
)
?
4'd3
:
(
SVRPkjTp
==
4'h7
)
?
4'd3
:
(
SVRPkjTp
==
4'h8
)
?
4'd7
:
(
SVRPkjTp
==
4'ha
)
?
4'd3
:
(
SVRPkjTp
==
4'hb
)
?
4'd7
:
4'd0
;
reg
[
3
:
0
]
SVRFuQLl
;
wire
[
1
:
0
]
SVRpkVSf
=
(
SVRFuQLl
==
4'd0
)
?
2'b00
:
(
SVRFuQLl
==
SVRYwUQz
)
?
2'b11
:
2'b01
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRFuQLl
<=
4'h0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRFuQLl
<=
4'bxxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRFuQLl
<=
4'h0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRpkVSf
==
2'b00
)
&&
SVRAyqoD
)
===
1'bx
)
SVRFuQLl
<=
4'bxxxx
;
`endif
else
if
(
(
SVRpkVSf
==
2'b00
)
&&
SVRAyqoD
)
SVRFuQLl
<=
4'd1
;
`ifdef SVRxoxPL 
else
if
(
(
SVRpkVSf
==
2'b01
)
===
1'bx
)
SVRFuQLl
<=
4'bxxxx
;
`endif
else
if
(
SVRpkVSf
==
2'b01
)
SVRFuQLl
<=
SVRFuQLl
+
4'd1
;
`ifdef SVRxoxPL 
else
if
(
(
SVRpkVSf
==
2'b10
)
===
1'bx
)
SVRFuQLl
<=
4'bxxxx
;
`endif
else
if
(
SVRpkVSf
==
2'b10
)
SVRFuQLl
<=
4'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRpkVSf
==
2'b11
)
===
1'bx
)
SVRFuQLl
<=
4'bxxxx
;
`endif
else
if
(
SVRpkVSf
==
2'b11
)
SVRFuQLl
<=
{
3'd0
,
SVRAyqoD
}
;
assign
SVRzfEzF
=
(
SVRYwUQz
==
4'd1
)
?
1'b1
:
(
SVRFuQLl
==
4'd0
)
?
1'b1
:
(
SVRFuQLl
==
SVRYwUQz
)
?
1'b1
:
1'b0
;
wire
[
15
:
0
]
SVRtyTOT
;
assign
SVRtyTOT
=
(
(
SVRPkjTp
==
4'h0
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
16'h0000
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
14'h0000
,
SVRMcPMP
[
7
:
6
]
}
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
14'b00_0000_0000_0000
,
SVRMcPMP
[
15
:
14
]
}
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
14'b00_0000_0000_0000
,
SVRMcPMP
[
23
:
22
]
}
:
(
SVRPkjTp
==
4'h1
)
?
{
14'b00_0000_0000_0000
,
SVRMcPMP
[
31
:
30
]
}
:
(
(
SVRPkjTp
==
4'h2
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
4'h0
,
SVRMcPMP
[
4
:
1
]
,
4'h0
,
SVRMcPMP
[
10
:
7
]
}
:
(
(
SVRPkjTp
==
4'h3
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
3'b000
,
SVRMcPMP
[
4
:
0
]
,
3'b000
,
SVRMcPMP
[
10
:
6
]
}
:
(
(
SVRPkjTp
==
4'h4
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
3'b000
,
SVRMcPMP
[
4
:
0
]
,
2'b00
,
SVRMcPMP
[
10
:
5
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
2'b00
,
SVRMcPMP
[
5
:
0
]
,
2'b00
,
SVRMcPMP
[
11
:
6
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
2'b00
,
SVRMcPMP
[
23
:
18
]
,
2'b00
,
SVRMcPMP
[
29
:
24
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
2'b00
,
SVRMcPMP
[
41
:
36
]
,
2'b00
,
SVRMcPMP
[
47
:
42
]
}
:
(
SVRPkjTp
==
4'h5
)
?
{
2'b00
,
SVRMcPMP
[
59
:
54
]
,
2'b00
,
SVRMcPMP
[
65
:
60
]
}
:
(
(
SVRPkjTp
==
4'h6
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
SVRMcPMP
[
7
:
0
]
,
SVRMcPMP
[
15
:
8
]
}
:
(
(
SVRPkjTp
==
4'h7
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
16'h0000
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
16'h0000
:
(
(
SVRPkjTp
==
4'ha
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
12'h000
,
SVRMcPMP
[
7
:
4
]
}
:
(
SVRPkjTp
==
4'ha
)
?
{
12'h000
,
SVRMcPMP
[
15
:
12
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
10'b00_0000_0000
,
SVRMcPMP
[
7
:
2
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
10'b00_0000_0000
,
SVRMcPMP
[
15
:
10
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
10'b00_0000_0000
,
SVRMcPMP
[
23
:
18
]
}
:
(
SVRPkjTp
==
4'hb
)
?
{
10'b00_0000_0000
,
SVRMcPMP
[
31
:
26
]
}
:
16'h0000
;
wire
[
7
:
0
]
SVRvFSMN
;
assign
SVRvFSMN
=
(
(
SVRPkjTp
==
4'h0
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
SVRMcPMP
[
7
:
0
]
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
SVRMcPMP
[
5
:
0
]
,
SVRMcPMP
[
33
:
32
]
}
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
SVRMcPMP
[
13
:
8
]
,
SVRMcPMP
[
35
:
34
]
}
:
(
(
SVRPkjTp
==
4'h1
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
SVRMcPMP
[
21
:
16
]
,
SVRMcPMP
[
37
:
36
]
}
:
(
SVRPkjTp
==
4'h1
)
?
{
SVRMcPMP
[
29
:
24
]
,
SVRMcPMP
[
39
:
38
]
}
:
(
(
SVRPkjTp
==
4'h2
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
4'h0
,
SVRMcPMP
[
15
:
12
]
}
:
(
(
SVRPkjTp
==
4'h3
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
3'h0
,
SVRMcPMP
[
15
:
11
]
}
:
(
(
SVRPkjTp
==
4'h4
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
3'h0
,
SVRMcPMP
[
15
:
11
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
2'h0
,
SVRMcPMP
[
17
:
12
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
2'h0
,
SVRMcPMP
[
35
:
30
]
}
:
(
(
SVRPkjTp
==
4'h5
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
2'h0
,
SVRMcPMP
[
53
:
48
]
}
:
(
SVRPkjTp
==
4'h5
)
?
{
2'h0
,
SVRMcPMP
[
71
:
66
]
}
:
(
(
SVRPkjTp
==
4'h6
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
SVRMcPMP
[
23
:
16
]
:
(
(
SVRPkjTp
==
4'h7
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
2'h0
,
SVRMcPMP
[
5
:
0
]
}
:
(
(
SVRPkjTp
==
4'h7
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
2'h0
,
SVRMcPMP
[
11
:
6
]
}
:
(
(
SVRPkjTp
==
4'h7
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
2'h0
,
SVRMcPMP
[
17
:
12
]
}
:
(
SVRPkjTp
==
4'h7
)
?
{
2'h0
,
SVRMcPMP
[
23
:
18
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
1'h0
,
SVRMcPMP
[
6
:
0
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
1'h0
,
SVRMcPMP
[
13
:
7
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
1'h0
,
SVRMcPMP
[
20
:
14
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h4
)
)
?
{
1'h0
,
SVRMcPMP
[
27
:
21
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h5
)
)
?
{
1'h0
,
SVRMcPMP
[
34
:
28
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h6
)
)
?
{
1'h0
,
SVRMcPMP
[
41
:
35
]
}
:
(
(
SVRPkjTp
==
4'h8
)
&&
(
SVRFuQLl
==
4'h7
)
)
?
{
1'h0
,
SVRMcPMP
[
48
:
42
]
}
:
(
SVRPkjTp
==
4'h8
)
?
{
1'h0
,
SVRMcPMP
[
55
:
49
]
}
:
(
(
SVRPkjTp
==
4'h9
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
SVRMcPMP
[
5
:
0
]
,
SVRMcPMP
[
33
:
32
]
}
:
(
(
SVRPkjTp
==
4'h9
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
SVRMcPMP
[
13
:
8
]
,
SVRMcPMP
[
35
:
34
]
}
:
(
(
SVRPkjTp
==
4'h9
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
SVRMcPMP
[
21
:
16
]
,
SVRMcPMP
[
37
:
36
]
}
:
(
SVRPkjTp
==
4'h9
)
?
{
SVRMcPMP
[
29
:
24
]
,
SVRMcPMP
[
39
:
38
]
}
:
(
(
SVRPkjTp
==
4'ha
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
SVRMcPMP
[
3
:
0
]
,
SVRMcPMP
[
19
:
16
]
}
:
(
SVRPkjTp
==
4'ha
)
?
{
SVRMcPMP
[
11
:
8
]
,
SVRMcPMP
[
23
:
20
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h1
)
)
?
{
SVRMcPMP
[
1
:
0
]
,
SVRMcPMP
[
37
:
32
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h2
)
)
?
{
SVRMcPMP
[
9
:
8
]
,
SVRMcPMP
[
43
:
38
]
}
:
(
(
SVRPkjTp
==
4'hb
)
&&
(
SVRFuQLl
==
4'h3
)
)
?
{
SVRMcPMP
[
17
:
16
]
,
SVRMcPMP
[
49
:
44
]
}
:
(
SVRPkjTp
==
4'hb
)
?
{
SVRMcPMP
[
25
:
24
]
,
SVRMcPMP
[
55
:
50
]
}
:
8'h00
;
reg
[
23
:
0
]
SVRdlnUs
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRdlnUs
<=
24'h000000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRdlnUs
<=
24'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRdlnUs
<=
24'h000000
;
else
SVRdlnUs
<=
{
SVRtyTOT
,
SVRvFSMN
}
;
reg
SVRxgbpl
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRxgbpl
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRxgbpl
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRxgbpl
<=
1'b0
;
else
SVRxgbpl
<=
(
SVRFuQLl
!=
4'd0
)
?
1'b1
:
1'b0
;
assign
SVRVmcEw
=
SVRdlnUs
;
reg
[
1
:
0
]
SVRWiSLk
;
reg
[
1
:
0
]
SVRyeWsF
;
always
@
(
SVRWiSLk
or
SVRoAAnA
or
SVRWTOHZ
or
SVRFuQLl
)
case
(
SVRWiSLk
)
2'd0
:
if
(
~SVRoAAnA
)
SVRyeWsF
=
2'd0
;
else
SVRyeWsF
=
2'd1
;
2'd1
:
if
(
SVRoAAnA
)
SVRyeWsF
=
2'd1
;
else
SVRyeWsF
=
2'd2
;
2'd2
:
if
(
SVRWTOHZ
)
SVRyeWsF
=
2'd2
;
else
SVRyeWsF
=
2'd3
;
2'd3
:
if
(
SVRFuQLl
!=
4'd0
)
SVRyeWsF
=
2'd3
;
else
SVRyeWsF
=
2'd0
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRWiSLk
<=
2'd0
;
else
if
(
SVRzUTNy
==
1'b1
)
SVRWiSLk
<=
2'd0
;
else
SVRWiSLk
<=
SVRyeWsF
;
assign
SVRoQJOJ
=
(
SVRWiSLk
!=
2'd3
)
?
1'b0
:
(
SVRyeWsF
!=
2'd0
)
?
1'b0
:
1'b1
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRfZzHt
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRGpakE
,
SVRcbwXF
,
SVRsgfsB
,
SVRvwyBE
,
SVRPQEPZ
,
SVRGolNq
,
SVRCAbmZ
,
SVRhVrUr
,
SVRklMnp
,
SVRBaLYP
,
SVRnAsZu
,
SVRFfTGh
,
SVRMxYWr
,
SVRbwSIu
)
;
input
wire
fclk
;
input
wire
SVRJROZz
;
input
wire
SVRzUTNy
;
input
wire
[
15
:
0
]
SVRGpakE
;
input
wire
SVRcbwXF
;
input
wire
SVRsgfsB
;
input
wire
SVRvwyBE
;
output
SVRPQEPZ
;
output
SVRGolNq
;
output
SVRCAbmZ
;
output
[
15
:
0
]
SVRhVrUr
;
output
[
7
:
0
]
SVRklMnp
;
output
[
15
:
0
]
SVRBaLYP
;
output
SVRnAsZu
;
output
SVRFfTGh
;
output
SVRMxYWr
;
output
SVRbwSIu
;
reg
[
7
:
0
]
SVRqYvKE
;
reg
[
7
:
0
]
SVRuSGkG
;
reg
[
7
:
0
]
SVRkwqfq
;
reg
[
7
:
0
]
SVRflIci
;
reg
SVRPQEPZ
;
reg
SVRGolNq
;
reg
SVRCAbmZ
;
reg
SVRMxYWr
;
wire
SVROYMTu
;
reg
[
1
:
0
]
SVRuzTwK
;
reg
[
1
:
0
]
SVRWFSdJ
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRWFSdJ
<=
2'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRWFSdJ
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
)
SVRWFSdJ
<=
2'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRWFSdJ
==
2'd3
)
===
1'bx
)
SVRWFSdJ
<=
2'bxx
;
`endif
else
if
(
SVRWFSdJ
==
2'd3
)
SVRWFSdJ
<=
2'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRsgfsB
==
1'd1
)
===
1'bx
)
SVRWFSdJ
<=
2'bxx
;
`endif
else
if
(
SVRsgfsB
==
1'd1
)
SVRWFSdJ
<=
2'd1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRWFSdJ
!=
3'd0
)
&&
(
SVRcbwXF
==
1'b1
)
)
===
1'bx
)
SVRWFSdJ
<=
2'bxx
;
`endif
else
if
(
(
SVRWFSdJ
!=
3'd0
)
&&
(
SVRcbwXF
==
1'b1
)
)
SVRWFSdJ
<=
SVRWFSdJ
+
2'd1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRMxYWr
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRMxYWr
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRMxYWr
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRMxYWr
==
1'b1
)
===
1'bx
)
SVRMxYWr
<=
1'bx
;
`endif
else
if
(
SVRMxYWr
==
1'b1
)
SVRMxYWr
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRcbwXF
==
1'b1
)
&&
(
SVRWFSdJ
==
2'd2
)
)
===
1'bx
)
SVRMxYWr
<=
1'bx
;
`endif
else
if
(
(
SVRcbwXF
==
1'b1
)
&&
(
SVRWFSdJ
==
2'd2
)
)
SVRMxYWr
<=
1'b1
;
else
SVRMxYWr
<=
1'b0
;
wire
[
7
:
0
]
SVRkjsuI
=
SVRGpakE
[
7
:
0
]
;
wire
[
7
:
0
]
SVRRXEci
=
SVRGpakE
[
15
:
8
]
;
wire
[
7
:
0
]
SVRVypbE
=
(
SVRvwyBE
==
1'b0
)
?
8'd0
:
(
SVRWFSdJ
==
2'd0
)
?
{
3'b000
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
3
]
^
SVRkjsuI
[
2
]
^
SVRkjsuI
[
1
]
,
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
3
]
^
SVRkjsuI
[
2
]
^
SVRkjsuI
[
0
]
,
SVRkjsuI
[
6
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
3
]
^
SVRkjsuI
[
1
]
^
SVRkjsuI
[
0
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
2
]
^
SVRkjsuI
[
1
]
^
SVRkjsuI
[
0
]
}
^
{
2'b00
,
SVRRXEci
[
7
]
^
SVRRXEci
[
6
]
^
SVRRXEci
[
5
]
^
SVRRXEci
[
4
]
^
SVRRXEci
[
3
]
^
SVRRXEci
[
2
]
,
SVRRXEci
[
1
]
^
SVRRXEci
[
0
]
,
SVRRXEci
[
7
]
^
SVRRXEci
[
6
]
^
SVRRXEci
[
5
]
^
SVRRXEci
[
1
]
^
SVRRXEci
[
0
]
,
SVRRXEci
[
7
]
^
SVRRXEci
[
4
]
^
SVRRXEci
[
3
]
^
SVRRXEci
[
1
]
,
SVRRXEci
[
6
]
^
SVRRXEci
[
4
]
^
SVRRXEci
[
2
]
^
SVRRXEci
[
0
]
,
SVRRXEci
[
5
]
^
SVRRXEci
[
3
]
^
SVRRXEci
[
2
]
}
:
(
SVRWFSdJ
==
2'd1
)
?
{
2'b00
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
3
]
^
SVRkjsuI
[
2
]
^
SVRkjsuI
[
1
]
^
SVRkjsuI
[
0
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
6
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
3
]
^
SVRkjsuI
[
2
]
^
SVRkjsuI
[
1
]
^
SVRkjsuI
[
0
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
3
]
,
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
2
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
1
]
,
SVRkjsuI
[
7
]
^
SVRkjsuI
[
6
]
^
SVRkjsuI
[
5
]
^
SVRkjsuI
[
4
]
^
SVRkjsuI
[
0
]
}
^
SVRRXEci
:
8'd0
;
wire
[
26
:
0
]
SVRxMHap
=
(
SVRvwyBE
==
1'b0
)
?
27'd0
:
(
SVRflIci
[
5
:
0
]
==
6'h00
)
?
27'h
4000000
:
(
SVRflIci
[
5
:
0
]
==
6'h07
)
?
27'h
2000001
:
(
SVRflIci
[
5
:
0
]
==
6'h0b
)
?
27'h
2000002
:
(
SVRflIci
[
5
:
0
]
==
6'h0d
)
?
27'h
2000004
:
(
SVRflIci
[
5
:
0
]
==
6'h0e
)
?
27'h
2000008
:
(
SVRflIci
[
5
:
0
]
==
6'h13
)
?
27'h
2000010
:
(
SVRflIci
[
5
:
0
]
==
6'h15
)
?
27'h
2000020
:
(
SVRflIci
[
5
:
0
]
==
6'h16
)
?
27'h
2000040
:
(
SVRflIci
[
5
:
0
]
==
6'h19
)
?
27'h
2000080
:
(
SVRflIci
[
5
:
0
]
==
6'h1a
)
?
27'h
2000100
:
(
SVRflIci
[
5
:
0
]
==
6'h1c
)
?
27'h
2000200
:
(
SVRflIci
[
5
:
0
]
==
6'h23
)
?
27'h
2000400
:
(
SVRflIci
[
5
:
0
]
==
6'h25
)
?
27'h
2000800
:
(
SVRflIci
[
5
:
0
]
==
6'h26
)
?
27'h
2001000
:
(
SVRflIci
[
5
:
0
]
==
6'h29
)
?
27'h
2002000
:
(
SVRflIci
[
5
:
0
]
==
6'h2a
)
?
27'h
2004000
:
(
SVRflIci
[
5
:
0
]
==
6'h2c
)
?
27'h
2008000
:
(
SVRflIci
[
5
:
0
]
==
6'h31
)
?
27'h
2010000
:
(
SVRflIci
[
5
:
0
]
==
6'h32
)
?
27'h
2020000
:
(
SVRflIci
[
5
:
0
]
==
6'h34
)
?
27'h
2040000
:
(
SVRflIci
[
5
:
0
]
==
6'h38
)
?
27'h
2080000
:
(
SVRflIci
[
5
:
0
]
==
6'h1f
)
?
27'h
2100000
:
(
SVRflIci
[
5
:
0
]
==
6'h2f
)
?
27'h
2200000
:
(
SVRflIci
[
5
:
0
]
==
6'h37
)
?
27'h
2400000
:
(
SVRflIci
[
5
:
0
]
==
6'h3b
)
?
27'h
2800000
:
(
SVRflIci
[
5
:
0
]
==
6'h01
)
?
27'h
2000000
:
(
SVRflIci
[
5
:
0
]
==
6'h02
)
?
27'h
2000000
:
(
SVRflIci
[
5
:
0
]
==
6'h04
)
?
27'h
2000000
:
(
SVRflIci
[
5
:
0
]
==
6'h08
)
?
27'h
2000000
:
(
SVRflIci
[
5
:
0
]
==
6'h10
)
?
27'h
2000000
:
(
SVRflIci
[
5
:
0
]
==
6'h20
)
?
27'h
2000000
:
27'h
1000000
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRqYvKE
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRqYvKE
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRqYvKE
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRWFSdJ
==
2'd0
)
&
(
SVRcbwXF
==
1'b1
)
)
===
1'bx
)
SVRqYvKE
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRWFSdJ
==
2'd0
)
&
(
SVRcbwXF
==
1'b1
)
)
SVRqYvKE
<=
SVRGpakE
[
7
:
0
]
;
reg
[
7
:
0
]
SVRklMnp
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRklMnp
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRklMnp
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRklMnp
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRWFSdJ
==
2'd2
)
===
1'bx
)
SVRklMnp
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRWFSdJ
==
2'd2
)
SVRklMnp
<=
SVRqYvKE
^
SVRxMHap
[
7
:
0
]
;
assign
SVROYMTu
=
(
SVRWFSdJ
==
2'd2
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRuzTwK
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRuzTwK
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
)
SVRuzTwK
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVROYMTu
==
1'b1
)
&&
(
SVRuzTwK
==
2'b00
)
)
===
1'bx
)
SVRuzTwK
<=
2'bxx
;
`endif
else
if
(
(
SVROYMTu
==
1'b1
)
&&
(
SVRuzTwK
==
2'b00
)
)
SVRuzTwK
<=
2'b01
;
`ifdef SVRxoxPL 
else
if
(
(
SVRuzTwK
==
2'b01
)
===
1'bx
)
SVRuzTwK
<=
2'bxx
;
`endif
else
if
(
SVRuzTwK
==
2'b01
)
SVRuzTwK
<=
2'b11
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVROYMTu
==
1'b0
)
&&
(
SVRuzTwK
[
0
]
==
1'b1
)
)
===
1'bx
)
SVRuzTwK
<=
2'bxx
;
`endif
else
if
(
(
SVROYMTu
==
1'b0
)
&&
(
SVRuzTwK
[
0
]
==
1'b1
)
)
SVRuzTwK
<=
2'b00
;
assign
SVRbwSIu
=
(
SVRuzTwK
==
2'b01
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRuSGkG
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRuSGkG
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRuSGkG
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRWFSdJ
==
2'd0
)
&
(
SVRcbwXF
==
1'b1
)
)
===
1'bx
)
SVRuSGkG
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRWFSdJ
==
2'd0
)
&
(
SVRcbwXF
==
1'b1
)
)
SVRuSGkG
<=
SVRGpakE
[
15
:
8
]
;
reg
[
7
:
0
]
SVRlTqAH
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRlTqAH
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRlTqAH
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRlTqAH
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRWFSdJ
==
2'd2
)
===
1'bx
)
SVRlTqAH
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRWFSdJ
==
2'd2
)
SVRlTqAH
<=
SVRuSGkG
^
SVRxMHap
[
15
:
8
]
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRkwqfq
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRkwqfq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRkwqfq
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRWFSdJ
==
2'd1
)
&
(
SVRcbwXF
==
1'b1
)
)
===
1'bx
)
SVRkwqfq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRWFSdJ
==
2'd1
)
&
(
SVRcbwXF
==
1'b1
)
)
SVRkwqfq
<=
SVRGpakE
[
7
:
0
]
;
reg
[
7
:
0
]
SVRFwiNq
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRFwiNq
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRFwiNq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRFwiNq
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRWFSdJ
==
2'd2
)
===
1'bx
)
SVRFwiNq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRWFSdJ
==
2'd2
)
SVRFwiNq
<=
SVRkwqfq
^
SVRxMHap
[
23
:
16
]
;
assign
SVRhVrUr
=
{
SVRFwiNq
,
SVRlTqAH
}
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRflIci
<=
8'haa
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRflIci
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
)
SVRflIci
<=
8'h00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRWFSdJ
==
3'd0
)
&
SVRcbwXF
)
===
1'bx
)
SVRflIci
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRWFSdJ
==
3'd0
)
&
SVRcbwXF
)
SVRflIci
<=
SVRVypbE
;
`ifdef SVRxoxPL 
else
if
(
(
SVRcbwXF
&
(
SVRWFSdJ
==
3'd1
)
)
===
1'bx
)
SVRflIci
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRcbwXF
&
(
SVRWFSdJ
==
3'd1
)
)
SVRflIci
<=
SVRflIci
^
SVRVypbE
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRPQEPZ
<=
1'b0
;
SVRGolNq
<=
1'b0
;
SVRCAbmZ
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
(
SVRzUTNy
==
1'b1
)
||
(
SVRvwyBE
==
1'b0
)
)
===
1'bx
)
begin
SVRPQEPZ
<=
1'bx
;
SVRGolNq
<=
1'bx
;
SVRCAbmZ
<=
1'bx
;
end
`endif
else
if
(
(
SVRzUTNy
==
1'b1
)
||
(
SVRvwyBE
==
1'b0
)
)
begin
SVRPQEPZ
<=
1'b0
;
SVRGolNq
<=
1'b0
;
SVRCAbmZ
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
(
SVRPQEPZ
==
1'b1
)
||
(
SVRGolNq
==
1'b1
)
||
(
SVRCAbmZ
==
1'b1
)
)
===
1'bx
)
begin
SVRPQEPZ
<=
1'bx
;
SVRGolNq
<=
1'bx
;
SVRCAbmZ
<=
1'bx
;
end
`endif
else
if
(
(
SVRPQEPZ
==
1'b1
)
||
(
SVRGolNq
==
1'b1
)
||
(
SVRCAbmZ
==
1'b1
)
)
begin
SVRPQEPZ
<=
1'b0
;
SVRGolNq
<=
1'b0
;
SVRCAbmZ
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRWFSdJ
==
2'd2
)
===
1'bx
)
begin
SVRPQEPZ
<=
1'bx
;
SVRGolNq
<=
1'bx
;
SVRCAbmZ
<=
1'bx
;
end
`endif
else
if
(
SVRWFSdJ
==
2'd2
)
begin
SVRPQEPZ
<=
SVRxMHap
[
26
]
;
SVRGolNq
<=
(
(
SVRxMHap
[
25
]
==
1'b1
)
|
(
SVRflIci
[
7
:
6
]
!=
2'b00
)
)
;
SVRCAbmZ
<=
SVRxMHap
[
24
]
;
end
reg
[
15
:
0
]
SVRBaLYP
;
reg
SVRnAsZu
;
reg
SVRFfTGh
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRBaLYP
<=
16'd0
;
SVRnAsZu
<=
1'b0
;
SVRFfTGh
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
begin
SVRBaLYP
<=
16'bxxxx_xxxx_xxxx_xxxx
;
SVRnAsZu
<=
1'bx
;
SVRFfTGh
<=
1'bx
;
end
`endif
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRBaLYP
<=
16'd0
;
SVRnAsZu
<=
1'b0
;
SVRFfTGh
<=
1'b0
;
end
else
begin
SVRBaLYP
<=
SVRGpakE
;
SVRnAsZu
<=
SVRcbwXF
;
SVRFfTGh
<=
SVRsgfsB
;
end
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRURDuX
(
fclk
,
pclk
,
SVRyEtuR
,
SVRWiNOI
,
SVRzUTNy
,
SVRrGCzn
,
SVRzMTVm
,
SVRehSHF
,
SVREusOH
,
SVRBdFMH
,
SVRmtjIy
,
SVRSCAjD
,
SVRklMnp
,
SVRjDxvg
,
SVREOLkD
,
SVRZmqEG
,
SVRBNOxF
,
SVRxmmsd
,
SVRbwSIu
,
SVRxZBBs
,
SVRXSjgA
,
SVRFoFlc
,
svr_cpu_int
)
;
input
fclk
;
input
pclk
;
input
SVRyEtuR
;
input
SVRWiNOI
;
input
SVRzUTNy
;
input
SVRrGCzn
;
input
SVRzMTVm
;
input
SVRehSHF
;
input
[
7
:
2
]
SVREusOH
;
input
[
7
:
2
]
SVRBdFMH
;
input
[
31
:
0
]
SVRmtjIy
;
input
SVRSCAjD
;
input
wire
[
7
:
0
]
SVRklMnp
;
input
wire
[
30
:
29
]
SVRjDxvg
;
input
wire
[
1
:
0
]
SVREOLkD
;
input
wire
[
30
:
28
]
SVRZmqEG
;
input
wire
[
30
:
29
]
SVRBNOxF
;
input
wire
[
15
:
0
]
SVRxmmsd
;
input
wire
SVRbwSIu
;
output
[
7
:
0
]
SVRxZBBs
;
output
[
31
:
0
]
SVRXSjgA
;
output
SVRFoFlc
;
output
svr_cpu_int
;
reg
[
7
:
0
]
SVRAyDvb
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRAyDvb
<=
8'hf8
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVREusOH
,
2'b00
}
==
`SVRmEdoF
)
)
===
1'bx
)
SVRAyDvb
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVREusOH
,
2'b00
}
==
`SVRmEdoF
)
)
SVRAyDvb
<=
SVRmtjIy
[
7
:
0
]
;
reg
[
7
:
0
]
SVRzFkDR
;
reg
[
7
:
0
]
SVRYibHm
;
reg
[
15
:
0
]
SVRzEAqG
;
wire
SVRyiJah
=
(
SVRbwSIu
==
1'b0
)
?
1'b0
:
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
?
1'b1
:
1'b0
;
wire
SVRyxNsU
=
(
SVRbwSIu
==
1'b0
)
?
1'b0
:
(
SVRklMnp
[
5
:
4
]
!=
2'b00
)
?
1'b1
:
1'b0
;
wire
SVRMLtjx
=
(
SVRjDxvg
[
29
]
==
1'b1
)
?
1'b1
:
(
SVREOLkD
[
1
:
0
]
==
2'b10
)
?
1'b1
:
(
SVRBNOxF
[
29
]
==
1'b1
)
?
1'b1
:
(
SVRZmqEG
[
28
]
==
1'b1
)
?
1'b1
:
1'b0
;
wire
SVRfMfxc
=
(
SVRBNOxF
[
30
]
==
1'b1
)
?
1'b1
:
(
SVRZmqEG
[
30
:
29
]
!=
2'b00
)
?
1'b1
:
(
SVREOLkD
[
1
:
0
]
==
2'b11
)
?
1'b1
:
(
SVRjDxvg
[
30
]
==
1'b1
)
?
1'b1
:
1'b0
;
wire
[
7
:
1
]
SVRcTClb
=
{
SVRyiJah
|
SVRzFkDR
[
7
]
,
SVRyxNsU
|
SVRzFkDR
[
6
]
,
1'b0
,
1'b0
,
1'b0
,
SVRMLtjx
|
SVRzFkDR
[
2
]
,
SVRfMfxc
|
SVRzFkDR
[
1
]
}
;
reg
SVRBwOFa
,
SVRzeqir
;
always
@
(
posedge
pclk
or
negedge
SVRWiNOI
)
if
(
~SVRWiNOI
)
SVRBwOFa
<=
1'b0
;
else
if
(
(
SVRzMTVm
==
1'b1
)
&&
(
SVRrGCzn
==
1'b1
)
&&
(
SVRSCAjD
==
1'b0
)
&&
(
{
SVRBdFMH
,
2'b00
}
==
`SVRgPbHP
)
)
SVRBwOFa
<=
1'b1
;
else
SVRBwOFa
<=
1'b0
;
always
@
(
posedge
pclk
or
negedge
SVRWiNOI
)
if
(
~SVRWiNOI
)
SVRzeqir
<=
1'b0
;
else
if
(
(
SVRzMTVm
==
1'b1
)
&&
(
SVRrGCzn
==
1'b1
)
&&
(
SVRSCAjD
==
1'b0
)
&&
(
{
SVRBdFMH
,
2'b00
}
==
`SVRPNWIl
)
)
SVRzeqir
<=
1'b1
;
else
SVRzeqir
<=
1'b0
;
wire
SVRmciEI
,
SVRgbepR
;
SVRPTXzm
SVRUWYmG
(
pclk
,
fclk
,
SVRBwOFa
,
SVRmciEI
)
;
SVRPTXzm
SVRJrVYG
(
pclk
,
fclk
,
SVRzeqir
,
SVRgbepR
)
;
reg
SVRdCTrH
,
SVRnHsBh
;
always
@
(
posedge
fclk
)
begin
SVRdCTrH
<=
SVRmciEI
;
SVRnHsBh
<=
SVRgbepR
;
end
wire
SVRSjfGu
=
(
SVRmciEI
&
(
~SVRdCTrH
)
)
;
wire
SVRWEcqK
=
(
SVRgbepR
&
(
~SVRnHsBh
)
)
;
wire
SVRFoFlc
=
SVRSjfGu
|
SVRWEcqK
;
reg
[
1
:
0
]
SVRKixaj
;
wire
SVRsElAe
=
(
SVRehSHF
==
1'b0
)
?
1'b0
:
(
{
SVREusOH
,
2'b00
}
==
`SVRgPbHP
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRKixaj
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRKixaj
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
)
SVRKixaj
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRsElAe
==
1'b1
)
===
1'bx
)
SVRKixaj
<=
2'bxx
;
`endif
else
if
(
SVRsElAe
==
1'b1
)
SVRKixaj
<=
{
SVRmtjIy
[
0
]
,
1'b0
}
;
else
if
(
(
SVRSjfGu
==
1'b1
)
&&
(
SVRKixaj
[
1
]
==
1'b0
)
)
SVRKixaj
<=
2'b00
;
else
if
(
(
SVRWEcqK
==
1'b1
)
&&
(
SVRKixaj
[
1
]
==
1'b0
)
)
SVRKixaj
<=
2'b00
;
else
if
(
(
SVRSjfGu
==
1'b1
)
&&
(
SVRKixaj
[
1
]
==
1'b1
)
)
SVRKixaj
<=
2'b11
;
else
if
(
(
SVRWEcqK
==
1'b1
)
&&
(
SVRKixaj
[
1
]
==
1'b1
)
)
SVRKixaj
<=
2'b11
;
else
if
(
SVRKixaj
==
2'b11
)
SVRKixaj
<=
2'b00
;
else
if
(
(
SVRKixaj
!=
2'b10
)
&&
(
SVRcTClb
[
7
:
1
]
!=
SVRzFkDR
[
7
:
1
]
)
)
SVRKixaj
<=
SVRKixaj
+
2'b01
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
begin
SVRzFkDR
<=
8'd0
;
SVRYibHm
<=
8'd0
;
SVRzEAqG
<=
16'd0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
begin
SVRzFkDR
<=
8'bxxxx_xxxx
;
SVRYibHm
<=
8'bxxxx_xxxx
;
SVRzEAqG
<=
16'bxxxx_xxxx_xxxx_xxxx
;
end
`endif
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRzFkDR
<=
8'd0
;
SVRYibHm
<=
8'd0
;
SVRzEAqG
<=
16'd0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRsElAe
==
1'b1
)
===
1'bx
)
begin
SVRzFkDR
<=
8'bxxxx_xxxx
;
SVRYibHm
<=
8'bxxxx_xxxx
;
SVRzEAqG
<=
16'bxxxx_xxxx_xxxx_xxxx
;
end
`endif
else
if
(
SVRsElAe
==
1'b1
)
begin
SVRzFkDR
<=
SVRmtjIy
[
7
:
0
]
;
SVRYibHm
<=
SVRmtjIy
[
15
:
8
]
;
SVRzEAqG
<=
SVRmtjIy
[
31
:
16
]
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
begin
SVRzFkDR
<=
8'bxxxx_xxxx
;
SVRYibHm
<=
8'bxxxx_xxxx
;
SVRzEAqG
<=
16'bxxxx_xxxx_xxxx_xxxx
;
end
`endif
else
if
(
SVRFoFlc
)
begin
SVRzFkDR
<=
8'd0
;
SVRYibHm
<=
8'd0
;
SVRzEAqG
<=
16'd0
;
end
else
begin
SVRzFkDR
<=
(
{
SVRcTClb
[
7
:
1
]
,
SVRKixaj
[
1
]
}
&
~SVRAyDvb
)
;
SVRYibHm
<=
SVRklMnp
;
SVRzEAqG
<=
SVRxmmsd
;
end
reg
SVRvIBfT
;
always
@
(
posedge
fclk
or
negedge
SVRyEtuR
)
if
(
SVRyEtuR
==
1'b0
)
SVRvIBfT
<=
1'b0
;
else
SVRvIBfT
<=
|
SVRzFkDR
[
7
:
1
]
;
assign
svr_cpu_int
=
SVRvIBfT
;
assign
SVRxZBBs
=
SVRAyDvb
;
assign
SVRXSjgA
=
{
SVRzEAqG
,
SVRYibHm
,
SVRzFkDR
}
;
endmodule
module SVRPTXzm
(
fclk
,
SVRkRNCW
,
SVRnXiwb
,
SVRSrADr
)
;
input
fclk
,
SVRkRNCW
,
SVRnXiwb
;
output
SVRSrADr
;
reg
SVRFVtoY
;
reg
SVRPXjhz
,
SVRUYEDm
;
reg
SVRxzPog
,
SVRLMuhd
;
always
@
(
posedge
fclk
)
if
(
SVRnXiwb
)
SVRFVtoY
<=
1'b1
;
else
if
(
SVRLMuhd
)
SVRFVtoY
<=
1'b0
;
always
@
(
posedge
SVRkRNCW
)
SVRPXjhz
<=
SVRFVtoY
;
always
@
(
posedge
SVRkRNCW
)
SVRUYEDm
<=
SVRPXjhz
;
always
@
(
posedge
fclk
)
SVRxzPog
<=
SVRUYEDm
;
always
@
(
posedge
fclk
)
SVRLMuhd
<=
SVRxzPog
;
assign
SVRSrADr
=
SVRUYEDm
;
initial
begin
SVRFVtoY
=
1'b0
;
SVRPXjhz
=
1'b0
;
SVRUYEDm
=
1'b0
;
SVRxzPog
=
1'b0
;
SVRLMuhd
=
1'b0
;
end
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRFwWBn
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRLwmmN
,
SVRhzkfv
,
SVRuPKrP
,
SVRJsIJK
,
SVRnckQL
,
SVRsUANj
,
SVRvqjMV
`ifdef SVRCadQw 
,
SVRCqyoW
,
SVRDmFCK
,
SVRjFeTQ
,
SVRQiYom
`endif
`ifdef SVReFgJe 
,
SVRCpDrC
,
SVRwBALo
,
SVRLnNsH
,
SVRSGtJq
`endif
`ifdef SVRaBkbf 
,
SVRMgbtT
,
SVRIJfkz
,
SVRdLyxD
,
SVRNliEf
`endif
)
;
input
wire
fclk
;
input
wire
SVRJROZz
;
input
wire
SVRzUTNy
;
input
wire
SVRLwmmN
;
input
wire
[
7
:
0
]
SVRhzkfv
;
input
wire
SVRuPKrP
;
input
wire
SVRJsIJK
;
output
wire
[
15
:
0
]
SVRnckQL
;
output
wire
SVRsUANj
;
output
SVRvqjMV
;
`ifdef SVRCadQw 
input
SVRCqyoW
;
input
[
7
:
0
]
SVRDmFCK
;
input
SVRjFeTQ
;
input
SVRQiYom
;
`endif
`ifdef SVReFgJe 
input
SVRCpDrC
;
input
[
7
:
0
]
SVRwBALo
;
input
SVRLnNsH
;
input
SVRSGtJq
;
`endif
`ifdef SVRaBkbf 
input
SVRMgbtT
;
input
[
7
:
0
]
SVRIJfkz
;
input
SVRdLyxD
;
input
SVRNliEf
;
`endif
`ifndef SVRCadQw
wire
SVRCqyoW
=
1'b0
;
`endif
`ifndef SVReFgJe
wire
SVRCpDrC
=
1'b0
;
`endif
`ifndef SVRaBkbf
wire
SVRMgbtT
=
1'b0
;
`endif
reg
[
15
:
0
]
SVRLvATy
;
reg
SVRSkNwM
;
wire
SVRwFtlt
=
(
SVRJsIJK
==
1'b1
)
?
1'b1
:
`ifdef SVRCadQw 
(
(
SVRCqyoW
==
1'b1
)
&&
(
SVRQiYom
==
1'b1
)
)
?
1'b1
:
`endif
`ifdef SVReFgJe 
(
(
SVRCpDrC
==
1'b1
)
&&
(
SVRSGtJq
==
1'b1
)
)
?
1'b1
:
`endif
`ifdef SVRaBkbf 
(
(
SVRMgbtT
==
1'b1
)
&&
(
SVRNliEf
==
1'b1
)
)
?
1'b1
:
`endif
1'b0
;
wire
[
1
:
0
]
SVRLPJFj
,
SVRSURPe
;
wire
SVRwXVuc
,
SVRXRTcS
;
wire
[
7
:
0
]
SVRYVwbw
,
SVRlrhTB
;
wire
[
3
:
0
]
SVRFIDWN
=
{
SVRMgbtT
,
(
~SVRMgbtT
)
&
(
SVRCpDrC
)
,
(
~SVRMgbtT
)
&
(
~SVRCpDrC
)
&
(
SVRCqyoW
)
,
(
~SVRMgbtT
)
&
(
~SVRCpDrC
)
&
(
~SVRCqyoW
)
}
;
wire
SVRBKKQK
=
SVRzUTNy
;
SVRnssvS
SVRscfdN
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRvuYtK
(
SVRhzkfv
[
7
:
0
]
)
,
.SVRwdvcj
(
SVRuPKrP
)
,
.read
(
SVRwXVuc
)
,
.SVRhTMHu
(
SVRwFtlt
)
,
.SVRHYuWd
(
SVRYVwbw
[
7
:
0
]
)
,
.SVRehbgg
(
SVRLPJFj
[
1
:
0
]
)
)
;
`ifdef SVRCadQw 
SVRnssvS
SVRCDadd
(
.fclk
(
fclk
)
,
.SVRJROZz
(
SVRJROZz
)
,
.SVRzUTNy
(
SVRzUTNy
)
,
.SVRvuYtK
(
SVRDmFCK
[
7
:
0
]
)
,
.SVRwdvcj
(
SVRjFeTQ
)
,
.read
(
SVRXRTcS
)
,
.SVRhTMHu
(
SVRwFtlt
)
,
.SVRHYuWd
(
SVRlrhTB
[
7
:
0
]
)
,
.SVRehbgg
(
SVRSURPe
[
1
:
0
]
)
)
;
`endif
localparam
SVROoABb
=
2'b00
;
localparam
SVRuhNNA
=
2'b01
;
localparam
SVRKDTtn
=
2'b11
;
localparam
SVReIsCX
=
1'b0
;
localparam
SVRokFGp
=
1'b1
;
localparam
SVRhFpQh
=
2'b00
;
localparam
SVRPIDNU
=
2'b01
;
localparam
SVRGKkmO
=
2'b10
;
localparam
SVRqsfgu
=
2'b11
;
localparam
SVRuCyVa
=
2'b00
;
localparam
SVRkoMxa
=
2'b01
;
localparam
SVRfhTla
=
2'b10
;
localparam
SVROwsYq
=
2'd1
;
localparam
SVRuljzI
=
2'd2
;
localparam
SVRfakxn
=
2'd3
;
wire
SVRKFEmR
=
(
(
SVRuPKrP
==
1'b1
)
||
(
SVRLPJFj
==
SVROwsYq
)
||
(
SVRLPJFj
==
SVRuljzI
)
)
;
`ifdef SVRCadQw 
wire
SVRSppGv
=
(
(
SVRjFeTQ
==
1'b1
)
||
(
SVRSURPe
==
SVROwsYq
)
||
(
SVRSURPe
==
SVRuljzI
)
)
;
`endif
reg
[
1
:
0
]
SVRiBDIb
,
SVRENoRA
;
always
@
(
*
)
case
(
SVRiBDIb
)
SVROoABb
:
if
(
SVRzUTNy
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
~SVRFIDWN
[
0
]
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRwFtlt
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRKFEmR
)
SVRENoRA
=
SVRuhNNA
;
else
SVRENoRA
=
SVROoABb
;
SVRuhNNA
:
if
(
SVRzUTNy
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRwFtlt
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRKFEmR
)
SVRENoRA
=
SVRKDTtn
;
else
SVRENoRA
=
SVRuhNNA
;
SVRKDTtn
:
if
(
SVRzUTNy
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRwFtlt
==
1'b1
)
SVRENoRA
=
SVROoABb
;
else
if
(
SVRKFEmR
)
SVRENoRA
=
SVRuhNNA
;
else
if
(
~SVRKFEmR
)
SVRENoRA
=
SVROoABb
;
else
SVRENoRA
=
SVROoABb
;
default
:
SVRENoRA
=
SVROoABb
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRiBDIb
<=
SVROoABb
;
else
if
(
SVRBKKQK
==
1'b1
)
SVRiBDIb
<=
SVROoABb
;
else
if
(
SVRLwmmN
==
1'b1
)
SVRiBDIb
<=
SVROoABb
;
else
if
(
SVRwFtlt
)
SVRiBDIb
<=
SVROoABb
;
else
SVRiBDIb
<=
SVRENoRA
;
`ifdef SVRCadQw 
reg
SVRbndoE
,
SVRMzxZF
;
always
@
(
*
)
case
(
SVRbndoE
)
SVReIsCX
:
if
(
SVRzUTNy
==
1'b1
)
SVRMzxZF
=
SVReIsCX
;
else
if
(
~SVRFIDWN
[
1
]
)
SVRMzxZF
=
SVReIsCX
;
else
if
(
SVRwFtlt
==
1'b1
)
SVRMzxZF
=
SVReIsCX
;
else
if
(
SVRKFEmR
&
SVRSppGv
)
SVRMzxZF
=
SVRokFGp
;
else
SVRMzxZF
=
SVReIsCX
;
SVRokFGp
:
if
(
SVRzUTNy
==
1'b1
)
SVRMzxZF
=
SVReIsCX
;
else
if
(
SVRwFtlt
==
1'b1
)
SVRMzxZF
=
SVReIsCX
;
else
if
(
~SVRKFEmR
&
~SVRSppGv
)
SVRMzxZF
=
SVReIsCX
;
else
SVRMzxZF
=
SVRbndoE
;
default
:
SVRMzxZF
=
SVReIsCX
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRbndoE
<=
SVReIsCX
;
else
if
(
SVRBKKQK
==
1'b1
)
SVRbndoE
<=
SVReIsCX
;
else
if
(
SVRLwmmN
==
1'b1
)
SVRbndoE
<=
SVReIsCX
;
else
if
(
SVRwFtlt
)
SVRbndoE
<=
SVReIsCX
;
else
SVRbndoE
<=
SVRMzxZF
;
`endif
assign
SVRwXVuc
=
(
SVRKFEmR
==
1'b0
)
?
1'b0
:
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b000
)
&&
(
SVRKFEmR
==
1'b1
)
)
?
1'b1
:
`ifdef SVRCadQw 
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b001
)
&&
(
SVRKFEmR
==
1'b1
)
&&
(
SVRSppGv
==
1'b1
)
)
?
1'b1
:
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b001
)
?
1'b0
:
`endif
`ifdef SVReFgJe 
(
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b01
)
&&
(
SVRfGhSg
!=
SVRoJzou
)
&&
(
SVRoJzou
!=
SVRqsfgu
)
)
?
1'b1
:
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b01
)
?
1'b0
:
`endif
`ifdef SVRaBkbf 
(
(
SVRMgbtT
==
1'b1
)
&&
(
SVRTKIZA
!=
SVRfhTla
)
&&
(
SVRwsRzN
==
SVRfhTla
)
)
?
1'b1
:
(
(
SVRMgbtT
==
1'b1
)
&&
(
SVRTKIZA
!=
SVRuCyVa
)
&&
(
SVRwsRzN
==
SVRuCyVa
)
)
?
1'b1
:
`endif
1'b0
;
`ifdef SVRCadQw 
assign
SVRXRTcS
=
(
SVRCqyoW
==
1'b0
)
?
1'b0
:
(
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b00
)
&&
(
SVRKFEmR
==
1'b1
)
&&
(
SVRSppGv
==
1'b1
)
)
?
1'b1
:
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b00
)
?
1'b0
:
`ifdef SVReFgJe 
(
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b01
)
&&
(
SVRfGhSg
!=
SVRoJzou
)
&&
(
SVRoJzou
!=
SVRGKkmO
)
)
?
1'b1
:
(
{
SVRMgbtT
,
SVRCpDrC
}
==
2'b01
)
?
1'b0
:
`endif
`ifdef SVRaBkbf 
(
(
SVRMgbtT
==
1'b1
)
&&
(
SVRTKIZA
!=
SVRfhTla
)
&&
(
SVRwsRzN
==
SVRfhTla
)
)
?
1'b1
:
(
(
SVRMgbtT
==
1'b1
)
&&
(
SVRTKIZA
!=
SVRuCyVa
)
&&
(
SVRwsRzN
==
SVRuCyVa
)
)
?
1'b1
:
`endif
1'b0
;
`endif
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRLvATy
<=
16'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRLvATy
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRLvATy
<=
16'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b000
)
&&
(
SVRENoRA
==
SVRuhNNA
)
&&
(
SVRwXVuc
==
1'b1
)
)
===
1'bx
)
SVRLvATy
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b000
)
&&
(
SVRENoRA
==
SVRuhNNA
)
&&
(
SVRwXVuc
==
1'b1
)
)
SVRLvATy
<=
{
8'd0
,
SVRYVwbw
}
;
`ifdef SVRxoxPL 
else
if
(
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b000
)
&&
(
SVRENoRA
==
SVRKDTtn
)
)
===
1'bx
)
SVRLvATy
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
{
SVRMgbtT
,
SVRCpDrC
,
SVRCqyoW
}
==
3'b000
)
&&
(
SVRENoRA
==
SVRKDTtn
)
)
SVRLvATy
<=
{
SVRYVwbw
,
SVRLvATy
[
7
:
0
]
}
;
`ifdef SVRCadQw 
`ifdef SVRxoxPL 
else
if
(
(
(
SVRMzxZF
==
SVRokFGp
)
)
===
1'bx
)
SVRLvATy
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRMzxZF
==
SVRokFGp
)
)
SVRLvATy
<=
{
SVRlrhTB
,
SVRYVwbw
}
;
`endif
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRSkNwM
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRENoRA
==
SVRuhNNA
)
)
===
1'bx
)
SVRSkNwM
<=
1'bx
;
`endif
else
if
(
(
SVRENoRA
==
SVRuhNNA
)
)
SVRSkNwM
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRwXVuc
==
1'b1
)
`ifdef SVRCadQw 
||
(
SVRXRTcS
==
1'b1
)
`endif
)
===
1'bx
)
SVRSkNwM
<=
1'bx
;
`endif
else
if
(
(
SVRwXVuc
==
1'b1
)
`ifdef SVRCadQw 
||
(
SVRXRTcS
==
1'b1
)
`endif
)
SVRSkNwM
<=
1'b1
;
else
SVRSkNwM
<=
1'b0
;
assign
SVRnckQL
=
SVRLvATy
;
assign
SVRsUANj
=
SVRSkNwM
;
reg
SVRxCrFk
,
SVRxHeiW
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRxCrFk
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
)
===
1'bx
)
SVRxCrFk
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
)
SVRxCrFk
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRxHeiW
==
1'b1
)
===
1'bx
)
SVRxCrFk
<=
1'bx
;
`endif
else
if
(
SVRxHeiW
==
1'b1
)
SVRxCrFk
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRLwmmN
==
1'b1
)
===
1'bx
)
SVRxCrFk
<=
1'bx
;
`endif
else
if
(
SVRLwmmN
==
1'b1
)
SVRxCrFk
<=
1'b1
;
wire
SVRvqjMV
=
(
SVRzUTNy
==
1'b1
)
?
1'b0
:
(
SVRxHeiW
==
1'b1
)
?
1'b0
:
(
(
SVRxCrFk
==
1'b1
)
&&
(
SVRsUANj
==
1'b1
)
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRxHeiW
<=
1'b0
;
else
SVRxHeiW
<=
SVRvqjMV
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRnssvS
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRvuYtK
,
SVRwdvcj
,
read
,
SVRhTMHu
,
SVRHYuWd
,
SVRehbgg
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRzUTNy
;
input
[
7
:
0
]
SVRvuYtK
;
input
SVRwdvcj
;
input
read
;
input
SVRhTMHu
;
output
[
7
:
0
]
SVRHYuWd
;
output
[
1
:
0
]
SVRehbgg
;
reg
[
7
:
0
]
SVRuSGkG
,
SVRkwqfq
;
reg
SVRfAYpj
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRfAYpj
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRfAYpj
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRfAYpj
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRhTMHu
)
===
1'bx
)
SVRfAYpj
<=
1'bx
;
`endif
else
if
(
SVRhTMHu
)
SVRfAYpj
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRwdvcj
==
1'b1
)
===
1'bx
)
SVRfAYpj
<=
1'bx
;
`endif
else
if
(
SVRwdvcj
==
1'b1
)
SVRfAYpj
<=
~SVRfAYpj
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRuSGkG
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRuSGkG
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRuSGkG
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRfAYpj
==
1'b0
)
&&
(
SVRwdvcj
==
1'b1
)
)
===
1'bx
)
SVRuSGkG
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRfAYpj
==
1'b0
)
&&
(
SVRwdvcj
==
1'b1
)
)
SVRuSGkG
<=
SVRvuYtK
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRkwqfq
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRkwqfq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRkwqfq
<=
8'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRfAYpj
==
1'b1
)
&&
(
SVRwdvcj
==
1'b1
)
)
===
1'bx
)
SVRkwqfq
<=
8'bxxxx_xxxx
;
`endif
else
if
(
(
SVRfAYpj
==
1'b1
)
&&
(
SVRwdvcj
==
1'b1
)
)
SVRkwqfq
<=
SVRvuYtK
;
parameter
SVRcnZHE
=
2'd0
;
parameter
SVROwsYq
=
2'd1
;
parameter
SVRuljzI
=
2'd2
;
parameter
SVRfakxn
=
2'd3
;
reg
[
1
:
0
]
SVRehbgg
,
SVRBGZqp
;
always
@
(
SVRehbgg
or
read
or
SVRwdvcj
)
case
(
SVRehbgg
)
SVRcnZHE
:
if
(
(
read
==
1'b0
)
&&
(
SVRwdvcj
==
1'b1
)
)
SVRBGZqp
=
SVROwsYq
;
else
if
(
(
read
==
1'b1
)
&&
(
SVRwdvcj
==
1'b0
)
)
SVRBGZqp
=
SVRfakxn
;
else
SVRBGZqp
=
SVRcnZHE
;
SVROwsYq
:
if
(
(
read
==
1'b0
)
&&
(
SVRwdvcj
==
1'b1
)
)
SVRBGZqp
=
SVRuljzI
;
else
if
(
(
read
==
1'b1
)
&&
(
SVRwdvcj
==
1'b0
)
)
SVRBGZqp
=
SVRcnZHE
;
else
SVRBGZqp
=
SVROwsYq
;
SVRuljzI
:
if
(
(
read
==
1'b0
)
&&
(
SVRwdvcj
==
1'b1
)
)
SVRBGZqp
=
SVRfakxn
;
else
if
(
(
read
==
1'b1
)
&&
(
SVRwdvcj
==
1'b0
)
)
SVRBGZqp
=
SVROwsYq
;
else
SVRBGZqp
=
SVRuljzI
;
default
:
SVRBGZqp
=
SVRfakxn
;
endcase
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRehbgg
<=
SVRcnZHE
;
else
if
(
SVRzUTNy
==
1'b1
)
SVRehbgg
<=
SVRcnZHE
;
else
if
(
SVRhTMHu
==
1'b1
)
SVRehbgg
<=
SVRcnZHE
;
else
SVRehbgg
<=
SVRBGZqp
;
assign
SVRHYuWd
=
(
SVRehbgg
==
SVRcnZHE
)
?
SVRvuYtK
:
(
(
SVRehbgg
==
SVROwsYq
)
&&
(
SVRfAYpj
==
1'b0
)
)
?
SVRkwqfq
:
(
(
SVRehbgg
==
SVROwsYq
)
&&
(
SVRfAYpj
==
1'b1
)
)
?
SVRuSGkG
:
(
(
SVRehbgg
==
SVRuljzI
)
&&
(
SVRfAYpj
==
1'b0
)
)
?
SVRuSGkG
:
SVRkwqfq
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
`define SVRiwKxv            6'b10_1010
`define SVRelSLK           6'b10_1011
`define SVRCfWss           6'b10_1100
module SVRalwrK
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRFoFlc
,
SVRehSHF
,
SVRyMsqX
,
SVRmtjIy
,
SVRUtdgF
,
SVRGolNq
,
SVRCAbmZ
,
SVRhVrUr
,
SVRFsZsI
,
SVRBCVbi
,
SVRnOXaE
,
SVRcbwXF
,
SVRsgfsB
,
SVRMxYWr
,
SVRgUyap
,
SVRpqIsy
,
SVRBaLYP
,
SVRnAsZu
,
SVRhirjM
,
SVRvwyBE
,
SVRpxeXJ
,
SVRHlCYR
,
SVRQfoZV
,
SVREOLkD
,
SVRBNOxF
,
SVRhWcSo
,
SVRxmmsd
,
SVRBcWQp
,
SVRDGtDt
,
SVRhnNgN
,
SVRGKeQn
,
SVRBAlYr
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRzUTNy
;
input
SVRFoFlc
;
input
SVRehSHF
;
input
[
7
:
2
]
SVRyMsqX
;
input
[
31
:
0
]
SVRmtjIy
;
input
[
16
:
5
]
SVRUtdgF
;
input
SVRGolNq
;
input
SVRCAbmZ
;
input
[
15
:
0
]
SVRhVrUr
;
input
[
7
:
0
]
SVRFsZsI
;
input
SVRBCVbi
;
input
[
15
:
0
]
SVRnOXaE
;
input
SVRcbwXF
;
input
SVRsgfsB
;
input
SVRMxYWr
;
output
[
7
:
0
]
SVRgUyap
;
output
reg
SVRpqIsy
;
output
[
15
:
0
]
SVRBaLYP
;
output
SVRnAsZu
;
output
SVRhirjM
;
input
SVRvwyBE
;
input
SVRpxeXJ
;
input
SVRHlCYR
;
input
SVRQfoZV
;
output
[
1
:
0
]
SVREOLkD
;
output
[
31
:
0
]
SVRBNOxF
;
output
SVRhWcSo
;
output
[
15
:
0
]
SVRxmmsd
;
output
wire
SVRBcWQp
;
output
SVRDGtDt
;
output
SVRhnNgN
;
output
[
5
:
0
]
SVRGKeQn
;
output
SVRBAlYr
;
wire
[
15
:
0
]
SVRwHBqh
=
SVRhVrUr
;
wire
SVRYgHNS
=
SVRpxeXJ
;
wire
SVRXJJAU
=
(
SVRYgHNS
==
1'b0
)
?
1'b0
:
1'b1
;
wire
SVRYRrnX
;
reg
[
31
:
0
]
SVRlPezP
;
reg
[
7
:
0
]
SVRgUyap
;
reg
[
15
:
0
]
SVRBaLYP
;
reg
SVRnAsZu
;
reg
SVRhirjM
;
reg
SVRFuCMU
;
reg
[
1
:
0
]
SVRpkotX
;
wire
SVRZfWeB
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRgUyap
<=
8'd0
;
SVRpqIsy
<=
1'b0
;
SVRBaLYP
<=
16'd0
;
SVRnAsZu
<=
1'd0
;
SVRhirjM
<=
1'd0
;
end
else
begin
SVRgUyap
<=
SVRFsZsI
;
SVRpqIsy
<=
SVRBCVbi
;
SVRBaLYP
<=
SVRnOXaE
;
SVRnAsZu
<=
(
SVRcbwXF
&
(
~SVRYRrnX
)
)
;
SVRhirjM
<=
SVRZfWeB
;
end
wire
[
5
:
0
]
SVRtYcCp
;
`ifdef SVRjzbOH 
wire
[
5
:
0
]
SVREMaUQ
=
SVRUtdgF
[
10
:
5
]
;
wire
[
5
:
0
]
SVRptaxv
=
SVRUtdgF
[
16
:
11
]
;
`ifdef SVRHjALk 
assign
SVRtYcCp
=
(
SVREMaUQ
==
6'd0
)
?
SVRFsZsI
[
5
:
0
]
:
(
SVRptaxv
==
6'd0
)
?
SVRFsZsI
[
5
:
0
]
:
(
SVRFsZsI
[
5
:
0
]
==
SVREMaUQ
)
?
SVRptaxv
:
SVRFsZsI
[
5
:
0
]
;
`else
assign
SVRtYcCp
=
(
SVREMaUQ
[
5
:
3
]
==
3'b010
)
?
SVRFsZsI
[
5
:
0
]
:
(
SVREMaUQ
[
5
:
4
]
==
2'b11
)
?
SVRFsZsI
[
5
:
0
]
:
(
(
SVRptaxv
!=
6'h22
)
&&
(
SVRptaxv
!=
6'h24
)
&&
(
SVRptaxv
!=
6'h2c
)
&&
(
SVRptaxv
!=
6'h2d
)
)
?
SVRFsZsI
[
5
:
0
]
:
(
SVRFsZsI
[
5
:
0
]
==
SVREMaUQ
)
?
SVRptaxv
:
SVRFsZsI
[
5
:
0
]
;
`endif
`else
assign
SVRtYcCp
=
SVRFsZsI
[
5
:
0
]
;
`endif
reg
[
5
:
0
]
SVRGKeQn
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRGKeQn
<=
6'd0
;
else
if
(
SVRBCVbi
)
SVRGKeQn
<=
SVRtYcCp
;
assign
SVRZfWeB
=
(
(
SVRFsZsI
[
5
:
4
]
!=
2'b00
)
&&
(
SVRMxYWr
==
1'b1
)
)
?
1'b1
:
1'b0
;
reg
[
14
:
0
]
SVRcYilW
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRcYilW
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRcYilW
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRcYilW
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRZfWeB
==
1'b1
)
===
1'bx
)
SVRcYilW
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRZfWeB
==
1'b1
)
SVRcYilW
<=
15'd1
;
`ifdef SVRxoxPL 
else
if
(
(
(
{
SVRcYilW
,
1'b0
}
<
(
SVRhVrUr
+
16'd2
)
)
&&
(
SVRcbwXF
==
1'b1
)
&&
(
SVRcYilW
!=
15'd0
)
)
===
1'bx
)
SVRcYilW
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
{
SVRcYilW
,
1'b0
}
<
(
SVRhVrUr
+
16'd2
)
)
&&
(
SVRcbwXF
==
1'b1
)
&&
(
SVRcYilW
!=
15'd0
)
)
SVRcYilW
<=
SVRcYilW
+
15'd1
;
`ifdef SVRxoxPL 
else
if
(
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRhVrUr
+
16'd2
)
)
===
1'bx
)
SVRcYilW
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRhVrUr
+
16'd2
)
)
SVRcYilW
<=
15'd0
;
reg
SVRnsaYo
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRnsaYo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRnsaYo
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRnsaYo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFsZsI
[
5
:
4
]
==
2'b00
)
===
1'bx
)
SVRnsaYo
<=
1'bx
;
`endif
else
if
(
SVRFsZsI
[
5
:
4
]
==
2'b00
)
SVRnsaYo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRnsaYo
==
1'b0
)
&&
(
{
SVRcYilW
,
1'b0
}
>=
SVRhVrUr
)
)
===
1'bx
)
SVRnsaYo
<=
1'bx
;
`endif
else
if
(
(
SVRnsaYo
==
1'b0
)
&&
(
{
SVRcYilW
,
1'b0
}
>=
SVRhVrUr
)
)
SVRnsaYo
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRnsaYo
==
1'b1
)
&&
(
SVRnAsZu
==
1'b1
)
)
===
1'bx
)
SVRnsaYo
<=
1'bx
;
`endif
else
if
(
(
SVRnsaYo
==
1'b1
)
&&
(
SVRnAsZu
==
1'b1
)
)
SVRnsaYo
<=
1'b0
;
wire
SVRscwrY
=
(
SVRFsZsI
[
5
:
4
]
==
2'b00
)
?
1'b0
:
(
(
{
SVRcYilW
,
1'b0
}
>=
SVRhVrUr
)
&&
(
SVRcbwXF
==
1'b1
)
&&
(
SVRcYilW
!=
15'd0
)
)
?
1'b1
:
1'b0
;
assign
SVRBcWQp
=
(
SVRFsZsI
[
5
:
4
]
==
2'b00
)
?
1'b0
:
(
SVRhVrUr
[
0
]
==
1'b0
)
?
1'b0
:
(
(
{
SVRcYilW
,
1'b0
}
>=
SVRhVrUr
)
&&
(
SVRnAsZu
==
1'b1
)
&&
(
SVRcYilW
!=
15'd0
)
)
?
1'b1
:
1'b0
;
reg
[
15
:
0
]
SVRxmmsd
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRxmmsd
<=
16'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRxmmsd
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRxmmsd
<=
16'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFuCMU
==
1'b1
)
===
1'bx
)
SVRxmmsd
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRFuCMU
==
1'b1
)
SVRxmmsd
<=
SVRhVrUr
;
reg
SVRvUgbq
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRvUgbq
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRvUgbq
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRvUgbq
<=
1'b0
;
else
if
(
SVRsgfsB
==
1'b1
)
SVRvUgbq
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRMxYWr
==
1'b1
)
&&
(
SVRZfWeB
==
1'b0
)
)
===
1'bx
)
SVRvUgbq
<=
1'bx
;
`endif
else
if
(
(
SVRMxYWr
==
1'b1
)
&&
(
SVRZfWeB
==
1'b0
)
)
SVRvUgbq
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFuCMU
==
1'b1
)
===
1'bx
)
SVRvUgbq
<=
1'bx
;
`endif
else
if
(
SVRFuCMU
==
1'b1
)
SVRvUgbq
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRXJJAU
==
1'b0
)
===
1'bx
)
SVRvUgbq
<=
1'bx
;
`endif
else
if
(
SVRXJJAU
==
1'b0
)
SVRvUgbq
<=
1'b0
;
reg
SVRkxDaI
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRkxDaI
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRkxDaI
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRkxDaI
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRyoryt
)
)
===
1'bx
)
SVRkxDaI
<=
1'bx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRyoryt
)
)
SVRkxDaI
<=
SVRmtjIy
[
8
]
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
SVRkxDaI
<=
1'bx
;
`endif
else
if
(
SVRFoFlc
)
SVRkxDaI
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRBCVbi
==
1'b1
)
&&
(
SVRFsZsI
[
5
:
0
]
==
6'd0
)
)
===
1'bx
)
SVRkxDaI
<=
1'bx
;
`endif
else
if
(
(
SVRBCVbi
==
1'b1
)
&&
(
SVRFsZsI
[
5
:
0
]
==
6'd0
)
)
SVRkxDaI
<=
SVRGolNq
;
reg
SVRoAAnA
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRoAAnA
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRoAAnA
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRoAAnA
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRZfWeB
==
1'b1
)
===
1'bx
)
SVRoAAnA
<=
1'bx
;
`endif
else
if
(
SVRZfWeB
==
1'b1
)
SVRoAAnA
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRhVrUr
+
16'd2
)
)
===
1'bx
)
SVRoAAnA
<=
1'bx
;
`endif
else
if
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRhVrUr
+
16'd2
)
)
SVRoAAnA
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRXJJAU
==
1'b0
)
===
1'bx
)
SVRoAAnA
<=
1'bx
;
`endif
else
if
(
SVRXJJAU
==
1'b0
)
SVRoAAnA
<=
1'b0
;
reg
SVRFLoar
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRFLoar
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRFLoar
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRFLoar
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRoAAnA
==
1'b1
)
&&
(
SVRXJJAU
==
1'b0
)
)
===
1'bx
)
SVRFLoar
<=
1'bx
;
`endif
else
if
(
(
SVRoAAnA
==
1'b1
)
&&
(
SVRXJJAU
==
1'b0
)
)
SVRFLoar
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRpkotX
==
2'b11
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
)
===
1'bx
)
SVRFLoar
<=
1'bx
;
`endif
else
if
(
(
SVRpkotX
==
2'b11
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
)
SVRFLoar
<=
1'b0
;
reg
SVRhWcSo
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRhWcSo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRhWcSo
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRhWcSo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRZfWeB
==
1'b1
)
===
1'bx
)
SVRhWcSo
<=
1'bx
;
`endif
else
if
(
SVRZfWeB
==
1'b1
)
SVRhWcSo
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
{
SVRcYilW
,
1'b0
}
>=
SVRwHBqh
)
===
1'bx
)
SVRhWcSo
<=
1'bx
;
`endif
else
if
(
{
SVRcYilW
,
1'b0
}
>=
SVRwHBqh
)
SVRhWcSo
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRXJJAU
==
1'b0
)
===
1'bx
)
SVRhWcSo
<=
1'bx
;
`endif
else
if
(
SVRXJJAU
==
1'b0
)
SVRhWcSo
<=
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRFuCMU
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRFuCMU
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRFuCMU
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRoAAnA
==
1'b1
)
&&
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRwHBqh
+
16'd2
)
)
)
===
1'bx
)
SVRFuCMU
<=
1'bx
;
`endif
else
if
(
(
SVRoAAnA
==
1'b1
)
&&
(
{
SVRcYilW
,
1'b0
}
>=
(
SVRwHBqh
+
16'd2
)
)
)
SVRFuCMU
<=
1'b1
;
else
SVRFuCMU
<=
1'b0
;
reg
[
15
:
0
]
SVRbmDsz
;
wire
[
15
:
0
]
SVRmzKBD
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRbmDsz
<=
16'h0000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRbmDsz
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRbmDsz
<=
16'h0000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRsgfsB
)
===
1'bx
)
SVRbmDsz
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRsgfsB
)
SVRbmDsz
<=
16'hffff
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRnAsZu
==
1'b1
)
&&
(
SVRoAAnA
==
1'b1
)
)
===
1'bx
)
SVRbmDsz
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRnAsZu
==
1'b1
)
&&
(
SVRoAAnA
==
1'b1
)
)
SVRbmDsz
<=
SVRmzKBD
;
wire
[
15
:
0
]
SVRGmSNo
=
(
SVRscwrY
==
1'b0
)
?
SVRnOXaE
:
(
SVRhVrUr
[
0
]
==
1'b0
)
?
SVRnOXaE
:
{
8'h00
,
SVRnOXaE
[
7
:
0
]
}
;
reg
[
15
:
0
]
SVRqgWth
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRqgWth
<=
16'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRqgWth
<=
16'bxxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRqgWth
<=
16'd0
;
else
SVRqgWth
<=
{
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
7
]
^
SVRGmSNo
[
15
-
3
]
,
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
6
]
^
SVRGmSNo
[
15
-
2
]
,
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
5
]
^
SVRGmSNo
[
15
-
1
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
7
]
^
SVRGmSNo
[
15
-
4
]
^
SVRGmSNo
[
15
-
0
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
6
]
,
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
5
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
4
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
7
]
^
SVRGmSNo
[
15
-
3
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
7
]
^
SVRGmSNo
[
15
-
6
]
^
SVRGmSNo
[
15
-
2
]
,
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
6
]
^
SVRGmSNo
[
15
-
5
]
^
SVRGmSNo
[
15
-
1
]
,
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
5
]
^
SVRGmSNo
[
15
-
4
]
^
SVRGmSNo
[
15
-
0
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
4
]
,
SVRGmSNo
[
15
-
15
]
^
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
7
]
^
SVRGmSNo
[
15
-
3
]
,
SVRGmSNo
[
15
-
14
]
^
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
10
]
^
SVRGmSNo
[
15
-
6
]
^
SVRGmSNo
[
15
-
2
]
,
SVRGmSNo
[
15
-
13
]
^
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
9
]
^
SVRGmSNo
[
15
-
5
]
^
SVRGmSNo
[
15
-
1
]
,
SVRGmSNo
[
15
-
12
]
^
SVRGmSNo
[
15
-
11
]
^
SVRGmSNo
[
15
-
8
]
^
SVRGmSNo
[
15
-
4
]
^
SVRGmSNo
[
15
-
0
]
}
;
assign
SVRmzKBD
[
0
]
=
SVRqgWth
[
0
]
^
SVRbmDsz
[
0
]
^
SVRbmDsz
[
4
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
12
]
;
assign
SVRmzKBD
[
1
]
=
SVRqgWth
[
1
]
^
SVRbmDsz
[
1
]
^
SVRbmDsz
[
5
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
13
]
;
assign
SVRmzKBD
[
2
]
=
SVRqgWth
[
2
]
^
SVRbmDsz
[
2
]
^
SVRbmDsz
[
6
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
13
]
^
SVRbmDsz
[
14
]
;
assign
SVRmzKBD
[
3
]
=
SVRqgWth
[
3
]
^
SVRbmDsz
[
3
]
^
SVRbmDsz
[
7
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
14
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
4
]
=
SVRqgWth
[
4
]
^
SVRbmDsz
[
4
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
5
]
=
SVRqgWth
[
5
]
^
SVRbmDsz
[
0
]
^
SVRbmDsz
[
4
]
^
SVRbmDsz
[
5
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
13
]
;
assign
SVRmzKBD
[
6
]
=
SVRqgWth
[
6
]
^
SVRbmDsz
[
1
]
^
SVRbmDsz
[
5
]
^
SVRbmDsz
[
6
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
13
]
^
SVRbmDsz
[
14
]
;
assign
SVRmzKBD
[
7
]
=
SVRqgWth
[
7
]
^
SVRbmDsz
[
2
]
^
SVRbmDsz
[
6
]
^
SVRbmDsz
[
7
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
13
]
^
SVRbmDsz
[
14
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
8
]
=
SVRqgWth
[
8
]
^
SVRbmDsz
[
3
]
^
SVRbmDsz
[
7
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
14
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
9
]
=
SVRqgWth
[
9
]
^
SVRbmDsz
[
4
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
12
]
^
SVRbmDsz
[
13
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
10
]
=
SVRqgWth
[
10
]
^
SVRbmDsz
[
5
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
13
]
^
SVRbmDsz
[
14
]
;
assign
SVRmzKBD
[
11
]
=
SVRqgWth
[
11
]
^
SVRbmDsz
[
6
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
11
]
^
SVRbmDsz
[
14
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
12
]
=
SVRqgWth
[
12
]
^
SVRbmDsz
[
0
]
^
SVRbmDsz
[
4
]
^
SVRbmDsz
[
7
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
15
]
;
assign
SVRmzKBD
[
13
]
=
SVRqgWth
[
13
]
^
SVRbmDsz
[
1
]
^
SVRbmDsz
[
5
]
^
SVRbmDsz
[
8
]
^
SVRbmDsz
[
9
]
;
assign
SVRmzKBD
[
14
]
=
SVRqgWth
[
14
]
^
SVRbmDsz
[
2
]
^
SVRbmDsz
[
6
]
^
SVRbmDsz
[
9
]
^
SVRbmDsz
[
10
]
;
assign
SVRmzKBD
[
15
]
=
SVRqgWth
[
15
]
^
SVRbmDsz
[
3
]
^
SVRbmDsz
[
7
]
^
SVRbmDsz
[
10
]
^
SVRbmDsz
[
11
]
;
wire
SVRuWtCu
=
(
SVRZfWeB
==
1'b1
)
?
1'b0
:
(
SVRmzKBD
==
16'h0000
)
?
1'b1
:
1'b0
;
reg
SVRBAlYr
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRBAlYr
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRnsaYo
==
1'b1
)
&&
(
SVRnAsZu
==
1'b1
)
&&
(
SVRuWtCu
!=
1'b1
)
)
===
1'bx
)
SVRBAlYr
<=
1'bx
;
`endif
else
if
(
(
SVRnsaYo
==
1'b1
)
&&
(
SVRnAsZu
==
1'b1
)
&&
(
SVRuWtCu
!=
1'b1
)
)
SVRBAlYr
<=
1'b1
;
`ifdef SVRxoxPL 
else
if
(
(
SVRsgfsB
==
1'b1
)
===
1'bx
)
SVRBAlYr
<=
1'bx
;
`endif
else
if
(
SVRsgfsB
==
1'b1
)
SVRBAlYr
<=
1'b0
;
reg
[
1
:
0
]
SVRkYjoK
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRkYjoK
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRWCIWM
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRWCIWM
)
)
SVRkYjoK
<=
SVRmtjIy
[
1
:
0
]
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRkYjoK
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
SVRFoFlc
)
SVRkYjoK
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRCAbmZ
==
1'b1
)
&&
(
SVRvwyBE
==
1'b1
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
(
SVRCAbmZ
==
1'b1
)
&&
(
SVRvwyBE
==
1'b1
)
)
SVRkYjoK
<=
2'b11
;
`ifdef SVRxoxPL 
else
if
(
(
SVRHlCYR
==
1'b1
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
SVRHlCYR
==
1'b1
)
SVRkYjoK
<=
2'b11
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRGolNq
==
1'b1
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
&&
(
SVRvwyBE
==
1'b1
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
(
SVRGolNq
==
1'b1
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
&&
(
SVRvwyBE
==
1'b1
)
)
SVRkYjoK
<=
2'b10
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRQfoZV
==
1'b1
)
&&
(
SVRhirjM
==
1'b1
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
(
SVRQfoZV
==
1'b1
)
&&
(
SVRhirjM
==
1'b1
)
)
SVRkYjoK
<=
2'b10
;
`ifdef SVRxoxPL 
else
if
(
(
(
(
SVRhirjM
==
1'b1
)
)
&&
(
SVRkYjoK
[
1
]
!=
1'b1
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
(
(
SVRhirjM
==
1'b1
)
)
&&
(
SVRkYjoK
[
1
]
!=
1'b1
)
)
SVRkYjoK
<=
2'b01
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRvUgbq
==
1'b0
)
&&
(
SVRkYjoK
!=
2'b11
)
)
===
1'bx
)
SVRkYjoK
<=
2'bxx
;
`endif
else
if
(
(
SVRvUgbq
==
1'b0
)
&&
(
SVRkYjoK
!=
2'b11
)
)
SVRkYjoK
<=
2'b00
;
reg
[
1
:
0
]
SVRfZehS
,
SVROsYVm
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRfZehS
<=
2'b00
;
SVROsYVm
<=
2'b00
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
begin
SVRfZehS
<=
2'bxx
;
SVROsYVm
<=
2'bxx
;
end
`endif
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRfZehS
<=
2'b00
;
SVROsYVm
<=
2'b00
;
end
else
begin
SVRfZehS
<=
SVRkYjoK
;
SVROsYVm
<=
SVRfZehS
;
end
assign
SVRYRrnX
=
~SVRvUgbq
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRpkotX
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRpkotX
<=
2'bxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRpkotX
<=
2'b00
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRvUgbq
==
1'b1
)
&&
(
SVRpkotX
==
2'b00
)
)
===
1'bx
)
SVRpkotX
<=
2'bxx
;
`endif
else
if
(
(
SVRvUgbq
==
1'b1
)
&&
(
SVRpkotX
==
2'b00
)
)
SVRpkotX
<=
2'b01
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRvUgbq
==
1'b0
)
&&
(
SVRpkotX
==
2'b01
)
)
===
1'bx
)
SVRpkotX
<=
2'bxx
;
`endif
else
if
(
(
SVRvUgbq
==
1'b0
)
&&
(
SVRpkotX
==
2'b01
)
)
SVRpkotX
<=
2'b10
;
`ifdef SVRxoxPL 
else
if
(
(
SVRpkotX
==
2'b10
)
===
1'bx
)
SVRpkotX
<=
2'bxx
;
`endif
else
if
(
SVRpkotX
==
2'b10
)
SVRpkotX
<=
2'b11
;
`ifdef SVRxoxPL 
else
if
(
(
SVRpkotX
==
2'b11
)
===
1'bx
)
SVRpkotX
<=
2'bxx
;
`endif
else
if
(
SVRpkotX
==
2'b11
)
SVRpkotX
<=
2'b00
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRlPezP
<=
32'h00000000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRlPezP
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRlPezP
<=
32'h00000000
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRyoryt
)
)
===
1'bx
)
SVRlPezP
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRyoryt
)
)
SVRlPezP
<=
SVRmtjIy
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
SVRlPezP
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRFoFlc
)
SVRlPezP
<=
32'h00000000
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRpkotX
==
2'b11
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
)
===
1'bx
)
SVRlPezP
<=
32'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRpkotX
==
2'b11
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
)
SVRlPezP
<=
{
(
~SVROsYVm
[
1
]
&
SVROsYVm
[
0
]
&
~
SVRBAlYr
&
~
(
SVRFsZsI
[
5
:
3
]
==
3'b111
)
&
~SVRFLoar
)
,
(
(
SVROsYVm
==
2'b11
)
|
(
SVRFsZsI
[
5
:
3
]
==
3'b111
)
|
SVRBAlYr
|
SVRFLoar
)
,
(
(
SVROsYVm
==
2'b10
)
|
(
SVRkxDaI
==
1'b1
)
)
,
SVRBAlYr
,
1'b0
,
SVRFLoar
,
1'b0
,
1'b0
,
1'b0
,
1'b0
,
1'b0
,
1'b0
,
11'd0
,
(
(
SVROsYVm
==
2'b10
)
|
(
SVRkxDaI
==
1'b1
)
)
,
SVRFsZsI
}
;
assign
SVREOLkD
=
SVRkYjoK
;
assign
SVRBNOxF
=
SVRlPezP
;
assign
SVRDGtDt
=
(
(
SVRpkotX
==
2'b11
)
&&
(
SVRFsZsI
[
5
:
3
]
!=
3'b000
)
)
?
1'b1
:
1'b0
;
assign
SVRhnNgN
=
(
(
SVRHlCYR
==
1'b1
)
&&
(
SVRkYjoK
!=
2'b11
)
)
?
1'b1
:
(
(
SVRGolNq
==
1'b1
)
&&
(
SVRkYjoK
!=
2'b10
)
)
?
1'b1
:
(
SVRhirjM
==
1'b1
)
?
1'b1
:
1'b0
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRBAPNY
(
fclk
,
SVRJROZz
,
SVRFoFlc
,
SVRehSHF
,
SVRyMsqX
,
SVRmtjIy
,
SVRmqigi
,
SVRLljSa
,
SVRYgHNS
,
SVRopDmx
,
SVROEvJE
,
`ifdef SVRCadQw 
SVRCqyoW
,
SVRTAKyC
,
SVRUxrba
,
`endif
SVRnCFbF
,
SVRjDxvg
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRFoFlc
;
input
SVRehSHF
;
input
[
7
:
2
]
SVRyMsqX
;
input
[
28
:
15
]
SVRmtjIy
;
input
SVRmqigi
;
input
SVRLljSa
;
input
SVRYgHNS
;
input
SVRopDmx
;
input
SVROEvJE
;
`ifdef SVRCadQw 
input
SVRCqyoW
;
input
SVRTAKyC
;
input
SVRUxrba
;
`endif
input
SVRnCFbF
;
output
[
31
:
15
]
SVRjDxvg
;
wire
SVRCpDrC
=
1'b0
;
wire
SVRDhaoC
=
1'b0
;
wire
SVROdaho
=
1'b0
;
wire
SVRMgbtT
=
1'b0
;
wire
SVRUbAdH
=
1'b0
;
wire
SVRXaNBq
=
1'b0
;
reg
[
28
:
15
]
SVRKtpgZ
,
SVRSJhDz
;
wire
SVRiLZGD
=
(
SVRLljSa
&
(
(
SVRKtpgZ
[
21
]
|
SVRKtpgZ
[
22
]
|
SVRKtpgZ
[
23
]
|
SVRKtpgZ
[
24
]
|
SVRKtpgZ
[
25
]
|
SVRKtpgZ
[
26
]
|
SVRKtpgZ
[
27
]
|
SVRKtpgZ
[
28
]
)
)
)
;
wire
SVRQLVIF
=
(
(
SVRLljSa
|
SVRCqyoW
|
SVRCpDrC
|
SVRMgbtT
)
&
(
SVRKtpgZ
[
16
]
|
SVRKtpgZ
[
17
]
|
SVRKtpgZ
[
18
]
|
SVRKtpgZ
[
19
]
|
SVRKtpgZ
[
20
]
)
)
;
wire
SVRhMTJg
=
(
SVRLljSa
&
(
~SVRiLZGD
)
&
(
~SVRQLVIF
)
)
;
reg
SVRdTWrD
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRdTWrD
<=
1'b0
;
else
SVRdTWrD
<=
SVRYgHNS
;
wire
SVRNpuBf
=
(
SVRYgHNS
==
1'b0
)
?
1'b0
:
(
SVRdTWrD
==
1'b1
)
?
1'b0
:
1'b1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRKtpgZ
<=
14'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRSfrTz
)
)
===
1'bx
)
SVRKtpgZ
<=
14'bxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRSfrTz
)
)
SVRKtpgZ
<=
SVRmtjIy
[
28
:
15
]
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
SVRKtpgZ
<=
14'bxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRFoFlc
)
SVRKtpgZ
<=
14'd0
;
else
SVRKtpgZ
<=
SVRSJhDz
;
always
@
(
*
)
SVRSJhDz
=
{
14
{
~SVRNpuBf
}
}
&
(
SVRKtpgZ
|
{
4'd0
,
SVRUbAdH
,
SVRDhaoC
,
SVRTAKyC
,
SVRopDmx
,
(
SVRnCFbF
&
SVRmqigi
)
,
SVRXaNBq
,
SVROdaho
,
SVRUxrba
,
SVROEvJE
,
1'b0
}
)
;
assign
SVRjDxvg
[
31
:
15
]
=
{
SVRhMTJg
,
SVRQLVIF
,
SVRiLZGD
,
SVRKtpgZ
[
28
:
15
]
}
;
endmodule
`define SVRfbgGT 
`define SVRCadQw 
`define SVRAtxnc 
`define SVRNJLgb 
`define SVRfLOvR 
`define SVRCsUKV  270000000
`define SVRojxSX  0
`define SVRJyIko      8'h00
`define SVRDfNXx         8'h04
`define SVRawpRC       8'h08
`define SVRmEdoF 	    8'h28
`define SVRgPbHP 	    8'h24
`define SVRPNWIl  8'h30
`define SVRgnUJW   8'h40
`define SVRPZskp   8'h44
`define SVRgtFxy   8'h48
`define SVRDJPlM   8'h4C
`define SVRORUft   8'h50
`define SVRUvXCJ    8'h54
`define SVRXKyOr     8'h58
`define SVRKlIMZ     8'h5C
`define SVRSfrTz         8'h80
`define SVRWCIWM   8'h84
`define SVRyoryt      8'h88
`define SVRmHiMj    8'h90
`define SVRGqeTe 	8'hA0
`define SVRqiCwc 	    8'hA4
`define SVRieolb 	    8'hA8
`define SVRqVcyR 	    8'hAC
`define SVRUqxEm        8'hF8
`define SVRJBHhX            8'hF0
`define SVRRNQDy            8'hF4
`define SVRhnrhd 		8'hFC
`define SVRDGIDb          8'hE0
`define SVRoqROa          8'hE4
`define SVRtBRmr          8'hE8
//`define SVRJNvGI 			   32'h01146101
`define SVRHElWy 
module SVRsbAVU
(
fclk
,
SVRJROZz
,
SVRzUTNy
,
SVRFoFlc
,
SVRehSHF
,
SVRyMsqX
,
SVRDtpEP
,
SVROJhPU
,
SVREOLkD
,
SVRBNOxF
,
SVRklMnp
,
SVRbwSIu
,
SVRvwyBE
,
SVRPQEPZ
,
SVRGolNq
,
SVRCAbmZ
,
SVRZmqEG
,
SVRDGtDt
,
SVRhnNgN
)
;
input
fclk
;
input
SVRJROZz
;
input
SVRzUTNy
;
input
SVRFoFlc
;
input
SVRehSHF
;
input
[
7
:
2
]
SVRyMsqX
;
input
[
31
:
17
]
SVRDtpEP
;
input
[
7
:
0
]
SVROJhPU
;
input
[
1
:
0
]
SVREOLkD
;
input
[
30
:
29
]
SVRBNOxF
;
input
[
7
:
0
]
SVRklMnp
;
input
SVRbwSIu
;
input
SVRvwyBE
;
input
SVRPQEPZ
;
input
SVRGolNq
;
input
SVRCAbmZ
;
output
[
31
:
0
]
SVRZmqEG
;
input
SVRDGtDt
;
input
SVRhnNgN
;
reg
[
8
:
0
]
SVRqPfym
;
wire
SVRIUcmg
;
parameter
SVRDqxYT
=
2'b00
;
parameter
SVRoIlZw
=
2'b01
;
parameter
SVRhRFzL
=
2'b11
;
parameter
SVRPOlFj
=
2'b10
;
reg
SVRuUFPE
;
reg
SVRwQlnG
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRuUFPE
<=
1'b0
;
SVRwQlnG
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
begin
SVRuUFPE
<=
1'bx
;
SVRwQlnG
<=
1'bx
;
end
`endif
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRuUFPE
<=
1'b0
;
SVRwQlnG
<=
1'b0
;
end
else
begin
SVRuUFPE
<=
SVRDGtDt
;
SVRwQlnG
<=
SVRhnNgN
;
end
reg
[
1
:
0
]
SVRxObZG
;
reg
[
1
:
0
]
SVRxNWrh
;
reg
[
1
:
0
]
SVRXmuBu
;
reg
[
1
:
0
]
SVRKZfgB
;
reg
SVRSZcDN
;
reg
SVRitXGk
;
reg
[
1
:
0
]
SVREJyqf
;
reg
[
1
:
0
]
SVRblIAT
;
reg
[
1
:
0
]
SVRAfrNW
;
reg
[
1
:
0
]
SVRZvemP
;
reg
SVRleyyL
;
reg
SVRfcmMs
;
reg
SVRcbgtj
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRleyyL
<=
1'b0
;
SVRfcmMs
<=
1'b0
;
SVRcbgtj
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
begin
SVRleyyL
<=
1'bx
;
SVRfcmMs
<=
1'bx
;
SVRcbgtj
<=
1'bx
;
end
`endif
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRleyyL
<=
1'b0
;
SVRfcmMs
<=
1'b0
;
SVRcbgtj
<=
1'b0
;
end
`ifdef SVRxoxPL 
else
if
(
(
SVRvwyBE
==
1'b0
)
===
1'bx
)
begin
SVRleyyL
<=
1'bx
;
SVRfcmMs
<=
1'bx
;
SVRcbgtj
<=
1'bx
;
end
`endif
else
if
(
SVRvwyBE
==
1'b0
)
begin
SVRleyyL
<=
1'b1
;
SVRfcmMs
<=
1'b0
;
SVRcbgtj
<=
1'b0
;
end
else
begin
SVRleyyL
<=
SVRPQEPZ
;
SVRfcmMs
<=
SVRGolNq
;
SVRcbgtj
<=
SVRCAbmZ
;
end
wire
SVRBaDJE
=
(
SVRZmqEG
[
7
:
0
]
!=
8'h00
)
?
1'b1
:
1'b0
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRqPfym
<=
9'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRqPfym
<=
9'bx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRqPfym
<=
9'd0
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRbwSIu
==
1'b1
)
&&
(
SVRklMnp
[
5
:
4
]
==
2'b00
)
)
===
1'bx
)
SVRqPfym
<=
9'bx_xxxx_xxxx
;
`endif
else
if
(
(
SVRbwSIu
==
1'b1
)
&&
(
SVRklMnp
[
5
:
4
]
==
2'b00
)
)
SVRqPfym
<=
{
SVRGolNq
,
SVRklMnp
}
;
wire
SVRhwAOL
=
(
(
SVRklMnp
[
5
:
0
]
==
6'd0
)
&
(
SVRbwSIu
==
1'b1
)
)
;
wire
SVRnAOrp
=
(
(
SVRhwAOL
==
1'b1
)
&&
(
SVRleyyL
==
1'b1
)
)
;
wire
SVRsgqBY
=
(
(
(
SVRitXGk
==
1'b1
)
&&
(
SVRBNOxF
[
30
]
==
1'b0
)
)
||
SVRFoFlc
)
;
wire
SVRvWdgq
=
(
(
SVRBNOxF
[
30
]
==
1'b0
)
&&
(
SVRBNOxF
[
29
]
==
1'b1
)
)
;
wire
SVRwRxVY
=
(
(
(
SVREOLkD
==
2'b11
)
&&
(
SVRwQlnG
)
)
||
(
(
SVRBNOxF
[
30
]
==
1'b1
)
&&
(
SVRuUFPE
)
)
||
(
(
SVRBNOxF
[
29
]
==
1'b1
)
&&
(
SVRuUFPE
)
)
)
;
wire
SVRLVLxz
=
(
SVRhwAOL
==
1'b1
)
;
wire
SVReRoEd
=
(
(
(
SVREOLkD
==
2'b11
)
&&
(
SVRwQlnG
)
)
||
(
(
SVRBNOxF
[
30
]
==
1'b1
)
&&
(
SVRuUFPE
)
)
)
;
wire
SVRCvhPb
=
(
(
SVRhwAOL
==
1'b1
)
&&
(
SVRcbgtj
==
1'b1
)
)
;
wire
SVROKDUa
=
(
(
SVRhwAOL
==
1'b1
)
&&
(
SVRfcmMs
==
1'b1
)
)
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
begin
SVRxObZG
<=
SVRDqxYT
;
SVRxNWrh
<=
SVRDqxYT
;
SVRXmuBu
<=
SVRDqxYT
;
SVRKZfgB
<=
SVRDqxYT
;
end
else
if
(
SVRzUTNy
==
1'b1
)
begin
SVRxObZG
<=
SVRDqxYT
;
SVRxNWrh
<=
SVRDqxYT
;
SVRXmuBu
<=
SVRDqxYT
;
SVRKZfgB
<=
SVRDqxYT
;
end
else
if
(
SVRFoFlc
&
~SVRBaDJE
)
begin
SVRxObZG
<=
SVRDqxYT
;
SVRxNWrh
<=
SVRDqxYT
;
SVRXmuBu
<=
SVRDqxYT
;
SVRKZfgB
<=
SVRDqxYT
;
end
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRmHiMj
)
)
begin
SVRxObZG
<=
SVROJhPU
[
1
:
0
]
;
SVRxNWrh
<=
SVROJhPU
[
3
:
2
]
;
SVRXmuBu
<=
SVROJhPU
[
5
:
4
]
;
SVRKZfgB
<=
SVROJhPU
[
7
:
6
]
;
end
else
if
(
SVRFoFlc
==
1'b1
)
begin
SVRxObZG
<=
SVRDqxYT
;
SVRxNWrh
<=
SVRDqxYT
;
SVRXmuBu
<=
SVRDqxYT
;
SVRKZfgB
<=
SVRDqxYT
;
end
else
begin
SVRxObZG
<=
SVREJyqf
;
SVRxNWrh
<=
SVRblIAT
;
SVRXmuBu
<=
SVRAfrNW
;
SVRKZfgB
<=
SVRZvemP
;
end
wire
[
2
:
0
]
SVRGLKpr
=
{
1'b0
,
SVRklMnp
[
7
:
6
]
}
;
wire
[
2
:
0
]
SVRQsSHI
=
{
1'b0
,
SVRklMnp
[
7
:
6
]
}
;
always
@
(
*
)
case
(
SVRxObZG
)
(
SVRDqxYT
)
:
if
(
(
SVRGLKpr
==
3'd0
)
&&
(
SVRnAOrp
==
1'b1
)
)
SVREJyqf
=
SVRoIlZw
;
else
if
(
(
SVRGLKpr
==
3'd0
)
&&
(
SVROKDUa
==
1'b1
)
)
SVREJyqf
=
SVRPOlFj
;
else
if
(
SVRQsSHI
!=
3'd0
)
SVREJyqf
=
SVRDqxYT
;
else
SVREJyqf
=
SVRDqxYT
;
(
SVRoIlZw
)
:
if
(
(
SVRGLKpr
==
3'd0
)
&&
(
SVRsgqBY
==
'b1
)
)
SVREJyqf
=
SVRDqxYT
;
else
if
(
(
SVRGLKpr
==
3'd0
)
&&
(
SVRLVLxz
==
'b1
)
)
SVREJyqf
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd0
)
SVREJyqf
=
SVRoIlZw
;
else
if
(
SVRvWdgq
==
1'b1
)
SVREJyqf
=
SVRPOlFj
;
else
if
(
SVRwRxVY
==
1'b1
)
SVREJyqf
=
SVRhRFzL
;
else
SVREJyqf
=
SVRoIlZw
;
(
SVRPOlFj
)
:
if
(
(
SVRGLKpr
==
3'd0
)
&&
(
SVRCvhPb
==
1'b1
)
)
SVREJyqf
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd0
)
SVREJyqf
=
SVRPOlFj
;
else
if
(
SVReRoEd
==
1'b1
)
SVREJyqf
=
SVRhRFzL
;
else
if
(
SVRsgqBY
==
1'b1
)
SVREJyqf
=
SVRDqxYT
;
else
SVREJyqf
=
SVRPOlFj
;
(
SVRhRFzL
)
:
if
(
SVRsgqBY
==
1'b1
)
SVREJyqf
=
SVRDqxYT
;
else
SVREJyqf
=
SVRhRFzL
;
default
:
SVREJyqf
=
SVRDqxYT
;
endcase
always
@
(
*
)
case
(
SVRxNWrh
)
(
SVRDqxYT
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRnAOrp
==
1'b1
)
)
SVRblIAT
=
SVRoIlZw
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVROKDUa
==
1'b1
)
)
SVRblIAT
=
SVRPOlFj
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRblIAT
=
SVRDqxYT
;
else
SVRblIAT
=
SVRDqxYT
;
(
SVRoIlZw
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRsgqBY
==
'b1
)
)
SVRblIAT
=
SVRDqxYT
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRLVLxz
==
'b1
)
)
SVRblIAT
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRblIAT
=
SVRoIlZw
;
else
if
(
SVRvWdgq
==
1'b1
)
SVRblIAT
=
SVRPOlFj
;
else
if
(
SVRwRxVY
==
1'b1
)
SVRblIAT
=
SVRhRFzL
;
else
SVRblIAT
=
SVRoIlZw
;
(
SVRPOlFj
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRCvhPb
==
1'b1
)
)
SVRblIAT
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRblIAT
=
SVRPOlFj
;
else
if
(
SVReRoEd
==
1'b1
)
SVRblIAT
=
SVRhRFzL
;
else
if
(
SVRsgqBY
==
1'b1
)
SVRblIAT
=
SVRDqxYT
;
else
SVRblIAT
=
SVRPOlFj
;
(
SVRhRFzL
)
:
if
(
SVRsgqBY
==
1'b1
)
SVRblIAT
=
SVRDqxYT
;
else
SVRblIAT
=
SVRhRFzL
;
default
:
SVRblIAT
=
SVRDqxYT
;
endcase
always
@
(
*
)
case
(
SVRXmuBu
)
(
SVRDqxYT
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRnAOrp
==
1'b1
)
)
SVRAfrNW
=
SVRoIlZw
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVROKDUa
==
1'b1
)
)
SVRAfrNW
=
SVRPOlFj
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRAfrNW
=
SVRDqxYT
;
else
SVRAfrNW
=
SVRDqxYT
;
(
SVRoIlZw
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRsgqBY
==
'b1
)
)
SVRAfrNW
=
SVRDqxYT
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRLVLxz
==
'b1
)
)
SVRAfrNW
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRAfrNW
=
SVRoIlZw
;
else
if
(
SVRvWdgq
==
1'b1
)
SVRAfrNW
=
SVRPOlFj
;
else
if
(
SVRwRxVY
==
1'b1
)
SVRAfrNW
=
SVRhRFzL
;
else
SVRAfrNW
=
SVRoIlZw
;
(
SVRPOlFj
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRCvhPb
==
1'b1
)
)
SVRAfrNW
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRAfrNW
=
SVRPOlFj
;
else
if
(
SVReRoEd
==
1'b1
)
SVRAfrNW
=
SVRhRFzL
;
else
if
(
SVRsgqBY
==
1'b1
)
SVRAfrNW
=
SVRDqxYT
;
else
SVRAfrNW
=
SVRPOlFj
;
(
SVRhRFzL
)
:
if
(
SVRsgqBY
==
1'b1
)
SVRAfrNW
=
SVRDqxYT
;
else
SVRAfrNW
=
SVRhRFzL
;
default
:
SVRAfrNW
=
SVRDqxYT
;
endcase
always
@
(
*
)
case
(
SVRKZfgB
)
(
SVRDqxYT
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRnAOrp
==
1'b1
)
)
SVRZvemP
=
SVRoIlZw
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVROKDUa
==
1'b1
)
)
SVRZvemP
=
SVRPOlFj
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRZvemP
=
SVRDqxYT
;
else
SVRZvemP
=
SVRDqxYT
;
(
SVRoIlZw
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRsgqBY
==
'b1
)
)
SVRZvemP
=
SVRDqxYT
;
else
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRLVLxz
==
'b1
)
)
SVRZvemP
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRZvemP
=
SVRoIlZw
;
else
if
(
SVRvWdgq
==
1'b1
)
SVRZvemP
=
SVRPOlFj
;
else
if
(
SVRwRxVY
==
1'b1
)
SVRZvemP
=
SVRhRFzL
;
else
SVRZvemP
=
SVRoIlZw
;
(
SVRPOlFj
)
:
if
(
(
SVRGLKpr
==
3'd1
)
&&
(
SVRCvhPb
==
1'b1
)
)
SVRZvemP
=
SVRhRFzL
;
else
if
(
SVRQsSHI
!=
3'd1
)
SVRZvemP
=
SVRPOlFj
;
else
if
(
SVReRoEd
==
1'b1
)
SVRZvemP
=
SVRhRFzL
;
else
if
(
SVRsgqBY
==
1'b1
)
SVRZvemP
=
SVRDqxYT
;
else
SVRZvemP
=
SVRPOlFj
;
(
SVRhRFzL
)
:
if
(
SVRsgqBY
==
1'b1
)
SVRZvemP
=
SVRDqxYT
;
else
SVRZvemP
=
SVRhRFzL
;
default
:
SVRZvemP
=
SVRDqxYT
;
endcase
reg
[
14
:
0
]
SVRvjWqR
;
assign
SVRIUcmg
=
(
SVRbwSIu
&
(
SVRklMnp
[
5
:
0
]
==
6'd1
)
)
;
wire
[
1
:
0
]
SVRKeyIv
=
(
SVRGLKpr
==
3'd0
)
?
SVRxObZG
:
(
SVRGLKpr
==
3'd1
)
?
SVRxNWrh
:
(
SVRGLKpr
==
3'd2
)
?
SVRXmuBu
:
(
SVRGLKpr
==
3'd3
)
?
SVRKZfgB
:
SVRxObZG
;
wire
[
1
:
0
]
SVRscmRk
=
SVRKeyIv
;
wire
SVRvUboW
=
(
SVRscmRk
[
1
:
0
]
==
SVRDqxYT
)
?
1'b1
:
1'b0
;
wire
SVRkXahy
=
(
SVRscmRk
[
1
:
0
]
==
SVRDqxYT
)
?
1'b0
:
1'b1
;
wire
SVRRrWVC
=
(
SVRscmRk
==
SVRhRFzL
)
?
1'b1
:
1'b0
;
wire
SVRViYxO
=
(
SVRscmRk
==
SVRPOlFj
)
?
1'b1
:
(
SVRGolNq
==
1'b1
)
?
1'b1
:
1'b0
;
wire
SVRxeZlU
=
(
SVRscmRk
!=
SVRoIlZw
)
?
1'b0
:
(
SVRGolNq
==
1'b1
)
?
1'b0
:
1'b1
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRvjWqR
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRvjWqR
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRFoFlc
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRFoFlc
)
SVRvjWqR
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRmHiMj
)
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRehSHF
&
(
{
SVRyMsqX
,
2'b00
}
==
`SVRmHiMj
)
)
SVRvjWqR
<=
SVRDtpEP
[
31
:
17
]
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRFoFlc
==
1'b1
)
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRFoFlc
==
1'b1
)
)
SVRvjWqR
<=
15'd0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRitXGk
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
SVRitXGk
)
SVRvjWqR
<=
{
SVRxeZlU
,
SVRvUboW
,
SVRRrWVC
,
SVRViYxO
,
SVRGLKpr
,
8'd0
}
;
`ifdef SVRxoxPL 
else
if
(
(
(
SVRhwAOL
==
1'b1
)
&&
(
SVRkXahy
==
1'b1
)
)
===
1'bx
)
SVRvjWqR
<=
15'bxxx_xxxx_xxxx_xxxx
;
`endif
else
if
(
(
SVRhwAOL
==
1'b1
)
&&
(
SVRkXahy
==
1'b1
)
)
SVRvjWqR
<=
(
SVRvjWqR
&
15'b1111_0001_1111_111
)
|
15'b0100_0000_0000_000
|
{
4'b0000
,
SVRGLKpr
,
8'b0000_0000
}
;
assign
SVRZmqEG
=
{
SVRvjWqR
,
SVRqPfym
[
8
:
0
]
,
SVRKZfgB
,
SVRXmuBu
,
SVRxNWrh
,
SVRxObZG
}
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRSZcDN
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRSZcDN
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRSZcDN
<=
1'b0
;
else
SVRSZcDN
<=
SVRIUcmg
;
always
@
(
posedge
fclk
or
negedge
SVRJROZz
)
if
(
SVRJROZz
==
1'b0
)
SVRitXGk
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRzUTNy
==
1'b1
)
===
1'bx
)
SVRitXGk
<=
1'bx
;
`endif
else
if
(
SVRzUTNy
==
1'b1
)
SVRitXGk
<=
1'b0
;
`ifdef SVRxoxPL 
else
if
(
(
SVRIUcmg
&
~SVRSZcDN
)
===
1'bx
)
SVRitXGk
<=
1'bx
;
`endif
else
if
(
SVRIUcmg
&
~SVRSZcDN
)
SVRitXGk
<=
1'b1
;
else
SVRitXGk
<=
1'b0
;
endmodule
module SVRBSVNR
(
SVRgYYWK
,
SVRtCTAv
,
SVRpsVqj
)
;
input
SVRgYYWK
;
input
SVRpsVqj
;
output
SVRtCTAv
;
reg
SVRsiYun
;
reg
SVRtCTAv
;
initial
#
0
begin
SVRsiYun
=
1'b0
;
SVRtCTAv
=
1'b0
;
end
always
@
(
posedge
SVRpsVqj
)
begin
SVRsiYun
<=
SVRgYYWK
;
SVRtCTAv
<=
SVRsiYun
;
end
endmodule